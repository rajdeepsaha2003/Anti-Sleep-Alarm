PK   ���WHX(�  Q�     cirkitFile.json�\�۸�W�W��"�[ӻ��^��݅AITV8�����A�����k�a�=�GQyX������=��W�����ξ�zU-������7��4�D�b�,g_j�p]}����������.��Ԓ�R�q*���d��VqB-�In���,���o'�;ű3;Ǳ�>�\*�.X,4�1�Y+�&�6��-)YR07%N�Ǯp��8,b��%H�$h	�d�I��fI���1/x�<�c�����~�c��c;���\�I�L��L�i),х�i��Y��<q�K�v[�bMJ'Vf����)u�m�7a��"#�I��Z�2�x�bC��Y�Z#�xA�7]�}Jf�Q� 79Enr��K�MN���"79H~�N��P$�)�=Q=f!�����z�ǐ�gHԳq�M���C�-�k��Zb�����X�@���u=6�(h�����790�̙�h>��������{扦\�<�Zd17I���H/�,+%��8Ȁ� ��H�ub�j'���F������qĶ�U�i<�����F�EJ�f��B�HaA�� R��R���!E�%"E��à.xà���/	�_�d��D$�T�h�Dm��4�i �4�iSF���Ɗ�bĄA1c�i��R$	�ğ,�Y�@�D�0(f'Q=�8n���t��6�P�.��������M��{]h�~bD�L�Ĉ���q+�S���9�������\�qDOiݪ1�Ŧu�nj3G�ux)4�D
"E�"�HI�HQA��0��0�%a�K����0	�`�$�I�0(�aPL��0(�aPLà��A1�b�4�i�0(faP��aP� ��D18��K9�N��pZ��rrD�/%�.'g��ᥜ8��K9�]hZ�����K���fS��U��ѕ�Dߪڮfs��b沾e]�:�����C����75�w�TȈ6���u ��q�2�#]�s@hu1>hl�a	sR1�3�B
�nF�<��(��,�aʀS���~OC���Zm�_�G3�bȹ];%_�����Q`�Q^�ߵ*�f���gR�+����E��  ���Q^$ �k������
�D��W ,��K�x�����p�cS�j�X�|��,��8��
lit�,�b�)��!�9��W&�LH ��H~���X8��$�"�`!I��$�d��fG*�����mvB�]EY1,l)ڎbaK���XضL�������Ӷn��Hd/`��-���8eX��#8'a�\��Ygp����uK�v�fGGV2G�\��3�i��L��UM�܃˛0c�s´<aځ+�qcm�ho�?&ѓ���霓�����Nz��g�oQ�<��z��(�G{���SOJ<-����a��OO<��s�V�砞�z�9�砞�z�9��ho�V��<k 
�>�CrL���� �����@y� ��C�z��m<f�_�� ���2f�b<*�8JԙLo��~3�2��F��Y@�{A�[����E��W���{�p�ﾋD�q �qg�O��׉�&�so(�2��m~����o۔��趉��ض��������ĶI���I�p��糬�n旦���r9�W�Ư�J�)�\�E�M�I!ݴJKB9�K�<�lFg������fs[6~�GD�����Mcܳ������Me�`��a���K�]5u����0���o�D_�|��y;^�<��u�����~]��ɍ�J3_Y׸���jUes�����^W�u�qp�qo���ͺ��1���4�����i������1Qt�@��Q&�����k���q_Ƅ�Y�\���bK�R�ϋ��Fq�}�"��,�(��D˺rkg6�Eu��qO���v���qJ�|_�t��P�$��\�*�*��L֗�����ZB���%�P��N�HM��6z���C|�n��߶M���Ѡ:롇�0H6��a�>���(��`����a�>��4L���Z07�q.1�%ǹ�(�P�D�Xt�x�6%�-�vP<Jl�@;=�G	������V5��uQ-?���)�R�O�YǖsE��p���n=�tj��J6�ľ-�2ͬ <N�b1wF�sZ�Tg�4$�"�][J|��|��7�L��v�U��<��d���f�����,��v/y��0e�����/���q#	�j�	g�������[%�&�}B�q��X��`���s"V,%��۔�y7���.nڐ�����>d������HI���v�6<;R��_ (�M(�D��J���� �T9w��.�S�8���,WҔ�кgV@']���Ӕ�k�-~���!}|��A2��|"{S��/�]p��~0��`����^�OEX"�i�H"]X�"��n�Ձ��.���%!%g��aIa�w�}LB�y�0ȱ(�q�6%�w"��Ym�ֿ�n�$����1K%} yW/M�$.\��xtgᝫr�-�R��f=aE�"e� q�
�����eb)r��&]��NāΊm !���Gˮ1��?�@���Kt��ܫ��S�ٽ��a������fҭ]Q� �ǹйզ�K��Rr��X�- ؤ=��{���PʴKy
N�Xm�^-�����ȥv[�N��.�I���V͝7�DL��wNw��U$������߻����C����������6��+��_��'����M����&��ٽW�&��8����X-�m���V�]GE�
J���|�R5'�p�=,�E��4w���777�?H����>��w�^]��7��1��9��Ty�IKǓ�d2L�N�����~8T�� +���s�{.���2:5LF���RP�g $���:�<C�W�!I:ba��2Ι�SЀ]4�#�L����ꝋ��4��d��:2 qw��>�[����A��K@h�j�|S�ϑdh�^F��D�n�a�1�aHn�N�*�U;#D?G�PV���%Oc�CEǢ/u�ll��+C.;��h�e�a��h��B��e�P���=���.M�@��F��t�[��V\���{[��5߇�h,~IAQ�!0�=�S�n9����:
�3�� g[�:
����$���(���jc��/��mD��7t�!�����!�F��1F�l$�n/�OFF|Qd��ət���S�o�n���C�=!�r�G�/<C;���.m���Dz��8u@��qѣ�v������_q��l���,}'�ӉAĥ�>b|��l$��u�j>���`[Wf���<�W��?��`k3���������я�PK   l��WK��( � /   images/967be514-0483-4001-9c2f-29bd6a1b95c6.png�{�S].�]�Yww��	���_���%Hp��,$@ x�@� �y������nWMM��s��L��~��C}MBzBm-�1�#0� >��'ܞL�o��ƚ�M����l7��*�iDwP��c-K�.�uW�`�?���`����L�����C�s��M2��<�Le(���Y�ր�k�U��碊�Z�SO�?�R@��S�Y_
8�߮.��3�,-=Q~�ɍ!�6��y�|�������$��0����ﬂ��[�w�BQ�K�'?d����'��X:l��S
MV0��F��O�%)�����b���J'��?��O�8���013��?�;�g�x��_��LH
@l�d��R�
/�@6���,lS�]�t�~��da�ҳ�M�5�d=���]�/n�7Ń?�\���J��~���V:�{~�	 ��W�c� ;�᛹�[hc++�Z�����j]��3���3�����N����{h��ŀ����&��!�$d�=I�W�5�el7q���U���L�p����O��F�LI��p42~dr+??�0���L8�5�N����F@�4	�w4}(��w�.x��Kn���?kC���$b���Jr��4��߾�Y}�)�B���/T��̣�U륬8����P�S&�?w|��e)>Ӕ��홧�;�U���~sc�^F|b5�u��k��8E
˷�#0�/q2�UlX0�Z�nZ���3Q�	��2�.E�r�1�?$��S������0��`�&�d�xh� z$q `-k8j!C�ҷ���M�ӄ���BFj�A����}�v��hf�NM�JMm-hx�V�&~�v��&�96-9��}��9)�|RϞ&��y�2�V�g�x��i���0E����w������'��BO�[��2�9Iji��9e�Se�P��ƕ��fX�g�^]�C�ч����.d�ͅ�؟�7	7$�qu���I�YP�b�{�e||�Vtu�����cHγ�B��JaN����i=nE�M��L)X���Ϫ��Y�u{�Y��oU��N�6K	���u9�'��6��������n��ʮ�Е����]��鯅'_:��z`|�pׯ��.Lr/��������K�ы&���/%����)	��(hzl�+C��;�}fH� ����d��r_��E׏�W�4��?�
1�}W)����B�-Jzћ�Ҽ������_o9�f�P_��yʨ^�݋+���m��Y�G���3Cdh�3���l���WW;o5�*�Y+�ܺӳ)&��Q�s��vag������c�� Jk����
h�h�{j��Z
`����f������S"�d��_�8T:\�)��Єޤ;zw5;�!��x#���e`�Hp�o5-�Q�����̯1B���0�Hi�\$r��>c$[�d���_���0�j!�%�����-v���:#�(%�F(Pu(��\Ugg���;� ?�ӄ�B��[�"��Nc$]��,�U�{�	��^����I&�$�"a�+���R+����Z}_����sE]��*,0�Y9>��b_�[u/��➐��}���N@��9�<?`a���������3�DE#s:���6̂��j��j\�Ы��j���h��eY�z��m�P��9<����137��䚫"ڟ�]�2���Sx�6<	�'��ZY�
oX���F"������s�} Q�i� �%2�hv���N9)�_�y�ߨg�ҥg��)s��m�������^��9��^�0w�
@�����p�ge~b�8��s�t� ;���έ���"/�����k{5� ğ3�<�* ��/�\��o�7�V�{R����������uwpͫj�Iu}���K�@5�V�J)��'���e]/C9f��'�3�G�ƪ�j���}y+���N��F�����;�QL0�o�g��Ѭ�(J�	�͗���srt!�N����U�&0���>U�����l1�=�`-�`��M"����^�0�ǅ������t�Ŏ��7rY؞���O/:Q��� 0���+u�vݒg��ŭX�dWm��
ee��+�/�!j������f}y3�]��j;!��C��/�[���.�u��t����/W���|�	�Wz3S�oTf�b�@��%��U�Y38Н�����Ë~������ m×&ci�10���d�J��ާ��E!ɪq0F{6�r��LK3�J,f^+���A���9��������R�ӛG�o�~$vUܽק��X��]]]��זQv0u�4t����@��k�>?��Dԭy����uRPa��{\d�n��0�%
1r�������rçܼZs�q"t_4k�iߌ�ĩ�L^ESꁞ����j�O@X��%)��W9�V����O*�d��d�8�4Y���'�wbE2�? Om=p�P�h��?�!�s����ji���TP�@V��4G2�����r���t}u�N�c��vU�W�4��w�E�Z|
7;&(�A��nv�����[�A]�ٰ�>����l쁿j2r;�!"6O�:�$2�$t���ŏ=
��aa�*2)7`EZ��
Q�h�ؓU!�~����z8�pX����Vt�"�^Ѥ�X$�.|���4xC�����}nT]��W�����2� �W�A��|���ʣeh�5D�Aǀ�Vm Ϩ�N'�S�;��� X�oeIW�ߘ�Fs���Vd��NJ�$<�٤��7ς��p�8�����b���\�#9zl:�����GG�^{�6=����w!����\;�桇�)_̰ꂞ\h�z�g� �������yfQƱ;Z$��^�H"�� ��Rb������[*�����_�S������o^�Pd&Ff=ǡl��+�0�� �W�9	�\:�%�����%�3�n2پ�N<�@�l�Ι5�އkWbǷ88)�r~����u@Aդ��uZ�����W7��rj�;/L	s�� I��&\iG�Т>�i�ٻ�(�ʒS���W.�_��]��)9G}aBB0��ڒف__Q�ƈ�%�\�n��ZAV�.����ю��������BߓJ��$��X%l�&�"��{
]��A���s��q�A�θ�a��Ku��[�{qf���� #���#���A�|O�U��h�	+���<z��[ܡ�rV�2��b�"Ľ��Y������p��]
wz�ы��QW���0�]w�n�}��K��g���L'����W>����� uM��1�	����~�=�2�r0���Q%%!Ѷ3F�ܒ�<��|}F%��2�b����J��ސa�[C�����3�+�9���p��?ECNGw����f�����N����q��&�f��~I�}L�$t5Q'dP���Z�J�Xl�9��Ru��W,k
���A��
��T�O-�9�[ڜ��^^s�f>����E5��N��Bم����>����ͨ�l��(�@�Fh��Ռ���R-D%�����M����lg$�R �����l�dD{����� 1u�ʗ�/"*`��Dov)))��ma�\ꢸ�Z������"�愢~4��0⳨HQG�w(�p�x�\���m���bAnE���*k�̻Ϗ(��h�#`���\࢏j��T +���zs%��-��m��NO��C@�?�����e�t�S�������ف�}�k���� �thVk��^m�V��l���"�Z�'�S#�$��:.7I�l�55��_Q��ܣ�Pߩ�i� �Md'���&C�e�3<��(ͷb�W����0��?|�}����m�ky��m��b�Q��V��*��Y�����ۢ=���/	��  ���" '�.L�X.�3L��8���î�����8��k�OX/���-mӕ\?��_��>Z�FE�V-���n��&<�>�͍d��f�%拍��eZ8��@c&4��_�� |>a�#��߭%�O5�՘,1�w�[lV��~_\o��	���PM��^ҷt���5*U��g J�l��M�;�F���j5�Y���R<19������T=��V�ŷuG�(}�
_�S�(Y���&��|D��������%P���Y�w�<�Wc�8L:��eO�fXd�s/om�j����^�$�zz��a�7ڹ��C�./ڕ~�w���ۯd�C�����;WU6�ӕ�īmա̩F���7�*�;�K�ʶJ 6����fL��6�4����'r#x��g�8?3Y����Q�a�]j/3�e�&f>'twRK:����:���L��o��/�Q�@ ��@�n��s4<Y�(y�ٓ�op�'����ǵT/�����c.L�ig~����?	����L�����v+R���ob���BP`&�^���9�F��S,d��gn����%V)�M�sn�^O��gV~��`�'}����Z7fn�[������k�E��������]��ŗ܅|���|����l�c���ܤq/N+��9j��Qp�(��lu��1T�P=��vao���_3v�1��峊�bH��4��2�6�8�����$d�+M_a �4�ጸjt��R%z����5�.Qb�i=A��߷`(���1<l�ř�v�;�`�z|�
��Hb�~^��Pi�������b+��ӥ�#��[tj��Wjq��<�zVAG�l�F�T��ؘ�S�f���kf؏��T�o�V�3���[�;�H2�?z~6y�C�l���(�kK�%�S�ψ(V�{������y>�s�1�0�K3��X��/A%6�_M����ܪ$�Đ�`��N��ʙJ�����%�����X���"H�j��}�����������0��a�n��V-��'��5��G^�yP���8�Z����*�O��q=�q�ao�[R��{n/
R�]�}�F�غ^�N���⨳�F՝���j��#���a�s�$#������ݒ`\��0��d��.���q�a����l��&����߫��U�����-���L@��ya�j�_E��D�����95�p���
9L|�'�|'L@�FE�P���1�7�A5�zy>��O�$�F����Y.gOݎ�z�D�$�A�B�Z�$�U�M�xw�_��3����I���K���w�o���S�cI��˗/�ygd{�А���ڧb����&ΩH�!�#9������P���\��Z;EH����t�j�Rt�2;��J���9$��Q�i��g��!%�zӳ�bk#�߇���7�!0�@l�y�lm�j=��vf3"�q��E���!����,L@.���#��G6�9oq���\��м�[����@~"��	1ښ&8��[O.�O�'��8(��-��� 3���������J�+چ��-�|�G��E�[w��*����Y[��ϳ��\i�Dn��4��
�]���tb�/��Ķ��Հw�^��Y��i�,�RѦ���p�ZcL̨�|�љK2z��~��9$�v�pة���qu��21]��/��ӰR�?���`ր�K�,�%���š���*e��Zr0�'�V�gKAXWW�ܷј�T/c�\E�r�G'���Qa8���-߇�O��{�F�O>?L�W�����_�~pi:&����@Q!�F��b�`�O6�6@6p/��.C!�a-�mqqa���q����$)z��XI`V@�̕]�er�jo�R���
Q5��.�'�yHf&vǾ�c}Sj9�,#[��Qn�sO���=��_yy_�M�f�Lܟ?���`����v�4߸����_g�)ͪ�2.�" `���p��ل
$�.H�P������'�W�a���l\���:n��/��1�I0�M���	��N*�����}У���տ&���ʈ�i=*%B�*��׿��}�@:wڽ���fm�������%��s�Ԯp[H�̔�6�o�!�<S�Kil���@JHR�G�yJթ��������O0 ��5��[��W���B�z��c�1
lK���AW��!W�Qz��g��p8zJ{�\Wu�ڦڅ��^����x�>-�ro��>�DNM��=4
�R��̙=���g����9�aN�����>MF%_�bk�b���؀�o�L긴��-�>�3Ղ��@iG3)x���~$��f��2L��8 �}�:ɻ�*��7�[��s�]/�cvC���a�k)G������A`=�a$ީ�Faܓ�c��w:������qU��6��I�~)��;�=ǉbR�y�����\���%M�ʏ	���D3�G�T-0��ӓ��&�~���H1��< �-���Pң����դ6���+?B�Tݔ��
n
�{�(�SZheR��e�!g^t�F�Gu�-P��ػڵ���/�A�j�sf!M6/L�/yLs��7���S\c��$�E�\JrMHy
��]/Vxz����=��U��oR��괟��_^?�����U.����UW`4f�N�&9��sv#�]�Rx�%��b�������\U��"�B
`��7���]�`��+�����de�*��,����%Ӗ7���6
�Ϥ���
���y���VH��V���l���Nv��8�q���$>���k�V���M��I�ذ��ј6���[q�]7�����}C���T!B����H�1O�CK턱�zN���5��i��*���b��f�x(�Q,W����X;�F��Ǌ������B��5��|��gq��,�(��3E?�b�=�1+k��_�j�iXC��7�wN~1�RרD��$d�i��<+�I��ճ�����	��W��!.�q�ʚڀ� V�ܸ4����պ�GX��Y���D�#�����~uM梵vǑ�I\�̐(�d�v�V���5]��$���;�m��$��+�{Ge��<f�o��=����*�O{�Bl��|1DȞ��y?�cb��M~�R��J���o �.+Cw�r������M_��8U���������B�nT�:�d��呥�M�H>4�r2�p]p�֍^X�(���7Y�ǯ 7�`�ѣ�m�S��N����'ZL�d�Àh�}]�v�,�J�FJ������GW�(8�-G�M�fw�	*��'�{�A�!��Cʦ�}Sod�ܵ|q���~�At�C~� u�ݗ��V��Y��=σ��GQ88�>�ܤZ��%�; ��HZ��2{q[�7?���aUk��2��q_�f+0�o���<��'Z$��[��r?P1[&���Q�����/��aY֘�9��ά#
M0ޣ�p�~2W$[,hӓn���ؚ�����M)�P��P���I��|3�+]DY+��8��Vy(6R�����E�=���G*@��nʤx"il��E>Ɛ7�ՑS�f��46��0|���+ri	�y�f�aK���j�fn��� �6)H�A�*�/�OcT驨�b��J�'vCb�Mo��!CC>5�dٗ���=����t��7������z�����(�P�D5�!v$+���ZAK��ր~CeN�[�#'����t��ęաA'��:I��^�����?�y��܆_.b�L�v7�6��酳+�<4$�d�7�M�hȠ������8��@Z<�^G�J��w�����+�� 7:��̄]��/yw��l3=��T���®�PE'�/�_�m�I<���\c�J/�Ŋ0^��`[�Of\ޡ�����m<!��#�x�&=�x���.;���\2dG*|��x��}��ܡQ���:[xm�B�i�&���p��O�P��K$ں|���8���yB}d&�<�а�5���)t�;���7���#�$Z��ҝ/<U~?����ϋ����^�m�O�[�ǆ(��;GU�=
�M��x:��".Nq����t�&�<��I�돏�X�.!�f����IL�gR�s���k(�12c�� 0�uVe.�OaJ�3
����L�h�����m@���6�/@E��5,E��8���=&9��?E	2x0d�c��6Z~O
uVD�״ʣ���,���Y��gu ��`c��.�0�)���#HB�i��������]�� N&�W���2��|��P��|���ڡ�0�ʭ.t���K�?2�v�ݵ�Y
�=r�(�O�5��6Pz�o�e����1Oc���g@�����k>�ֽ4�Z��Ic�y���?������Ƶ����^llt��f��\{T�|�s�%�4�x*:q�R �d����S��#=���0�X�W-4�PYA�a=џ�S�I$W�ʿ	MH���u8�r���g@�W�MG~H�9�W��� ,��7n�|���No(*6�./ԛ���Yq����4��g�z:�+�\��o�,�^8�l=��J��+`G��tA~�X��s6F�ZW�.GGO��ό����:E�S��>�.��<��]�'W\�L"��Ɔ����_���z�3��d��{����?�Y7��09��tM�`����;f�;��
��Gі1���H�e�\vr�~ޗ}�����������i��u3�>�=���?����0E)b��|z�<���u p�Eȩ��� �.�PM��B��b�]�����Ƶ�,W��K����7�JTP��/�������ߤ�a��nJ�9��ŋX�7[����Ԍ~씨^�ͥ:�vn�,sqŉ*��$�&��6J��3�PqGW[�=����n�=���"��1H�T�]�d��.�}�{珬�}i��G�Ha]q����w���̪upN��䕱�����x���f�����ݞ�j�,�>��v���w�~�z�7�!k��; ���L�t�����*�;��ij���65���<#�;v<��`%�zY�j�g���khKY:����P�A	"<���Š��pU�<~���q�<{�RJ�|�����W�F""��/��Hs�z�LWo���5i��H3�vU���`�� �=���y�"R�CD�p��D�,.�.��ď;!�{G�<��~�K� ����̗"�h�7·jjK��o��k�����������]�ڬ9����x��Y�GJ�,��	����o��m�  �.�n�{[�_�s�o8��ka�z�#"4@����g�7!�U��gVWY���-f
��9���<�p|�\�C�ߪe�_�vI���p�ly,�HdkX��LԄ�G����B=��65��F�/�X�����Xh]V�d��l�>��F���8ڨV�Hu��S�L=�4��ݖjj7w�{�R�`�Ģ^�Q9��ךT̴�K��������G> �_���y��ǪӺp��;,�+��1�ѩ���W�Z�7��t�� k�;J��NW�1�|^�'VjP���Ԫqx^��r8i���}ϼ2�s g�8/m�@�c�
7ˋ�@�L��q��`\�j�'Χ�P��㼁�m�AMN�.n�IB����1a`�<��qU6������|�<@-��<\� qsr2�V�gZ�h�;�4�o(X�tr��6WrY/�*3�tH:f���%xI4@e!�fnQˍuP��Y�.%����̺�?U?t�wl�1nJ|=�%���a±6T�v6�=��r��M'�����gч.&YY��i �1ŕq�}�7϶�4$��&��/r/a�R�4�)���P��R�(~~Y���aʏt�x���j��&��@����Z��� �� &�S��
.~d��E��9Kvr���'��Q�:G41*ō�C)^ �6���)���9	���GSY��ճ;TraM��Gţ�)y<����>�i8��v��|Y�D
��}��e�q~W�}]�nR���Αc�ʅ���xCQ1�ۊ��*�$�X-iy��b��WD�j�?IC��T~��m�E�c=�W���*5���$o���3�)�tс�\}&{f�{*?O�_�RV��~u:�H�M��#��T����:���Y��uX�>2��"�O��,q�]y��UM�ɚp��b���E�N#S����M�z;�
����̓��cδu:�F�m~�o��K�q�P0���P"<X��_�W�D�
�p�����[0x��/>�꧳����J�S#[��?��EPp�c�n�PUH^!t�S]=���� �*v�Վ���+��2'Rܢ�q[�э�[������s�-�R\�$3ד��f~���ǆ��h��&�O�����������0�L*x���C���f[��Y�+�Q�d�fю�^��w~ՙ~*U,!��ī&���`Љ�i�i��5a�^ S�!��w����2�B>��V��
�1v�b�#�����v�t�#���o�e������TWK��%C�!�?�_�Sc�,��#�ʷ&76GOb]&7ӚxY,�؋�oϋ����l
a=%}��3R`��Q�(W�ݯh�d���/�����AO��v��g�g��}u��"20G�b� I���L�],j������E�p��ΎK[��ӽ?�
�@����g��n~����Q�dV��z	=TN�Fo�7~��A����P��X� �䵯�_�����g�����5B���eqtb!܅�#X�U��:�q�[�=
�ldXe�gia��Ȯ�9�VM�Cb�j��p�Gy��ޅ���'�ޅd�6fZ��
 S��#a~�2n��J�h��]����^k�OD�%�kG�Ʀ{B���է�T��N"l|R�s5�dyڒ
B]o���+;��*LdNv�y\!q�1z�[����q7-4p<�*�w9�b�҇U�a��i�;X�� ��gm� �=K�1��J%�Ǎ<;I���\P���F�^�x\�a�Ff��ڴ�	� � ?�H�s.1g:��]��e]��LQ,�5_}���%�B�����;���"3�ϛC��j��h�����\�X�P�����0 Kx�`�p|��p�l*�bV75�>T�����!��R�2�/B+�Lv8Vn�;��_'Ŵ���߯�ⴿ$j����'��:f�L���˰�'�U�Ocj���BJ�a7ˋk���S�=��D�R��]½���a�D�ǧY���AS�Da�%����)H�xVk���S�]$IY6u������S����Ǜx��RQ~i8�-ҹ��C��^!��/rZ�r<4��=j��,�x��WKe|+�jb:R��EW=$☨���s3���U��v.B
n:f��� XV��61�๟:��=)I}��z���eP/N��g �3��9���������%8��h���iu�ڷ��r���5ׅ�4w���^_/��r��h�t	jٙaE&��3#%���*�F�p{/F>g5�}d�{ �c��"𕢜�U��6���Sm�B��m 	�� �t�8:)II���-F��t�w����J��B)��;��%&��s��獿�=���^�w@h槶��3ik�J�x�f�;B<%l�m�Vw1^/�}_{u���sI�>�����Fw��c,sl1����f�_u��:H:�ܥ�7��z\�5G�TJj��c��Ck�TE�ۂh����1�}�+p��Ǒ��*$���J��`�;�뗜�4G5��d�r�b��n��׮�S�~��kZ:���>īm
�ܪ�)-�*1��5�+��GA�\�7fA"��H��x�5��xx{%>v=����s-�|�¾����h�,�ǈ��g���THk�Z���N��w68����͢j�3x:txg=ofr�%�-�΅�q�Hw�
)D �[-c^��P�k�LMg�о
@��㫪���C�����l��I;w��I���R���C�� ��;��	ر[�'�H�)C@�����&�]H�ŋSv?���;�*Tb^{��n�����s��̣����>))�/#���z�hq~H��o����/^��f���|�v�fm��d҈�;#M�E�e:��v'�إ�P+��p"�s'y���|��R�X���O��;�?\(���P��T����^R&���
ӧ-�oY������"�����Gb�k��7g�q����DV^��]ƗO.�O��?}�}I�wQY�_8
��ݬb81]�w���b��h�@��uy���}�������_�O�K�D'/z�G��N¨���D1e�h����Ԡ�pi-l�k��0��Md�Q�L��`	�3(L[SI�8��^��=L{���������0�=� ��
r�m��Cfhf1Y�7���W�B�x�:U�N���n�)xu[��J/(�_��=%��� ��nG#��(uw�mf��)giT՘��^[t�Uf�S'���-C��>�3��l��Oa�G��8�����ݡ���U�Xē#^MNp۩�~��3�
|5]���b��a�*0;�u���Ҷ��N<�?+i��7���� �0
Y��Y����,li�����?t���֌����4�uzwb�r�8ֻ}�4�΃4zS����=�:⃆����������
�C�����]Dwo���N5������'��EZ��V��W��w1��d���1q��w��e��!y�2�}��Vj�U���;�p�}4!Z�l�*��ֱ��Ba���!�cYȊ���N��s	4ӟ�Fl|��r��/�ov��u�V��Fn�T��K%];�+�t:��n���z)TI8C(MU�����f"��6Y�r�.$	���,���s�+�͔D��`W����B	�ؔ�W��k�T �q�6���!��dޢ:gg>�t���M(��B���E��nV7�«��M��1�+���:�[Z����@�B{�"�W�-��2�;P0؏�8M�hCs�2��̲�]GF�������ī�Gk��ï����ۂ����<����K��s�x{�������`���M	����ܝ��Rכ-V�>O�@�6����u�ǘ��E4�}Rk�">�X&�^f�i���w{�	�B)��?�|��ț{�.Kߧt�������NW�{������}���ǳƥ`/G��5����=q��gyr�{O�<[1������;M�� ����{�^<}�����,�v�έ��Λ8��k���EՌ�ˬ��FG�����?%l���P����_�[[)��`u��,}E��)LX�j���`���sD���@f$�*8��T+�Q$y��Y�hCB��A���L�O�zvΡ�9T���̄���s���4��+;D"0�����G��捄�3�� 2�xebĦw���{u�[vఛQ�j� |tC��y"ߴ��6I�s�>3��.�Ǹ\�n��*{O'�Z�����9�|ʖ}5G�H,�6S���6���>O�P�����R���24X�!4��>~,�ǂ����d�\6+|Z�^{;�w���T�t�uuUw`�i=V����^��W�6�e1@��*�;q~X�L�`;��m��fe7�s�r�v�������y=�k�!
0��_��^�Z]G�X'���:��I������2�v�$:R�tgI�`9�u��\���bII����m�Y�Cw���/y�xYE�x5 �����xzCSS�X9}�`-9���L-S԰�Pe@6?��۔0n�9�l�ʛ~,DD`��]�+nL��f�)J^
��ٕå�c�V�w޴ 03��l�R�B������l|l/4�F|����(9^4��b�2�y�C���)v��w����|B۵�g�}�����!)	��Θo�<��4��T@&�\��F�+S��r�1��ڮP�Q���^ԃ�����,��={��iQ��MT�,���N)��4����K1K�ﭨc�k��if�%�]*I�nʆ�d���GW5\Œ��uWp�w|`�ZZ&���	�����s"0:�i3ޚ�/��������;�=��Q����P��cߋ�V}����\GQ��ϸ+&Õ�y�YD:�0-(M
���ؙ�4V;��Q�u&�|���s��Aq
�[����܅3��bI4��n���r����M�mL��+��888��� � (A���Q�:J��9g�Q�68��21:�����]*�,R5�>�h�)*�[b^��~n�4�;%�q��>�m���򨻠)L�
��m�[�s��"�z�zB����ǣ,"�8z������4>p�A�R�^5���AY9qp�8^�I���纄jXZXE+�����E�B�VQڤ��Y�[�=��<b��4�у83v~�+ϧ�CB�^��z?w�;Y0�+�fN�)8p����r���M<4��c���yp�{Ć3��ͦ
�)��������E eWd_��ĥ�q}���|�%�Ҧk����Gn�ऋ�M�`&h�+K��5-s�u];��U�c7j���9ꧽi�&dj�F.�<�)����?><׿�T��p�@MnBu�P���S�Kx|��`��"�"��I�j��:(u�;�z�gh����ow_��o�(d�\����ݸw0L�D�w's!0����h�]-6V=٤<��?b��@D^�+�w%��1%�?�!�����/4{)-�4
�$ls!�K	~��nWψG��?:�D�J��,��G�x��/彮t��$�;���i-�F�7����tT���{�[1d���(/h���4n,�[?��c�����N��͸�K�X�7&��tB�x����*�)���kN6�\QU�o� �LuB'�C�,�z(���P�l����wH����m"-�3��d#;�nNG
�e�<�u-��8�n���K5<u��<]&�HوF�-	oӇ
�}���WLW��Tx�d�e��V5!M&�K���<�c]����{~���f�D-�����/�d���(�����a�S��u^h9�+�W+����La���e;�� �ғBa|f[��OO��j��C��Ӄ%а���ݸׇ4�D��/_���s��Z�8%�M��?R��$8Zd<�g���H�>\�<|�51���s�@���ة���ܻV�ަ�$i�,@gug*?�48����!HMJ�����u��E�4l�;?p�o}I��t�ѩ�}����I�[B��׃`�D�ŕ���WP���vSlCWϚ�SRC7.�x߻��.�^��~������^D��/�G������i=�Vw�Vַ��y_9���63�vr	����7I��2(��gߧ&l%�M���(�����u�|��O�����a\���[A�ps�Z0���}�u��O�����IXr5��S��|8q��\�r*��B�\V���,G(;1@��{��S����(�FӦB�&çꢽ��\��:[s��u��Yn6z��Ա��r7aX�.�3���M��`IjZ/k�N��ȅ�ږ��Mv�l����y-?����H���}S<����H*8P�S���N�6�G#dI��dhO4���1���W�(GG�:��v�����c8��ܻ��p,W�k�{w_ud��kV}p�n��(����m�G��d�d��ܨN�)z&�eU���<Q̜į}�S-w^��i��oq�d���G��>��=\U����b5%����Ύ����e@�>��(��A�a���۷�̠��兟_�B� �OTgh�Jy��z�;��đ/��5���v��Igj+�6���11qV��i�g��,b̘y��4�cV �M�-N	n���4i	��f��ѿ�,T��(5��a�_?�՚�Bb�X��ܿ&��8{k�#�=�	�Y�/'&ɤ���ԎIM1��P���F�{�4�I��'`E�<a�4��UPX��wzX�.�sS��c�4�u�9f�h'r���hiA�Q3�%PZv;W�������pɈ�������W�����/@�KLe���:�\xa�iN ��o-�P-�MH��� Ն��my׶���Z�k�h�k_�B?Ƈ����4�\��s
ln�̅+���=4 ���K�(.G%\3~��;�V�����G�/.�Hj�Y�x�"N��c^ ��c���i��:0?�y��-���#���tgC�:��c�x�Xbq�;k\�Q�z�6�-��պ���ϴ̩?�R�r'������_Vl��1p���?�y�E�I�
��z��E�e����;e�.��;J��F*�̢g>��V!n�"d��5�/��?�LX�6E��O�8cR^D-��;9	9�b������zuCЫ�T����q��ǽ�4b���fe�ݍ��*Uo�A)N�'�|� p��w/F�Q��*�@WX��%� p���	��e�NZ@�&\���q�JZ��������d~����b�yl���Ў�2��j��I�
qg�=;�3�[�o=K'+��q���% =fG0�-��+�&�0��s�%RN1�/�\M��յ3ʅi(L����&
���;�2�����(ي�����!ԭ����1}�r��K鐡�R�����v{]��l�y�;?+�m�)RVG:�t�㏶m�J�z5r���M�sr
����,�[�O5�	��K��</��B_S��p'�f�lr��d�{� �@l���(cv���:��͛�_��������+�����n$Q�}m�⽉Z��vw�i�}L�;c�4���<fw�{�̓i���\�=W�
�=��0�R���E�<����wm=�����܁�c-���ԭ�y���Nn���	��#,7U<���cY����<��
�_lF`n����D���ē5��$F���G���`-���h&��"� ���2��OG��J���Ӥx�/E���*�/JKq�a���2�|���G���i<$/��T}�r.ɭ�,paSN$�2	���~OR��4� �y6�$0"�$X�G�ǎ�����Ξ�1�U�Fr�O��b�q[u�\&�bƒ⹅e=�o���.�6����k���~�o�nZ^ZV�2J��7z�\�Ik��noZ�/Dka~w�/�#eΫ�������G�����g��}ԛG�ys�Ə1������޽{&%�{;�8��{�y����6u��2��ܖ�c��N�n��_�tVz�H�2��l�y�un�L
 � >4�lB�0n=�V���cs����Di��EqI��	�Vd(yK@2�|�-��d����nH	��ɲ?A�C�LDt� U����al�/2 %�〬q�?���!�D�GVWу�a|"B���|���"��:7�.lQk��������9g"	a��R�W�?��8� �Y�1D�<��Tԣ��ˤ�`����b�{�`�%���]#D��X6�w>���%������(CHr����R>�j�Cr�)_{�|��DD��<oda~>�9s�o�}��t�����˶�dxN�²X��|����>}����A!"B4��&����?�Q���Mn��?_���=5�,Uf��^?�Y�U䭷�M?��[��w�NW�^��H���͗���}R3�EG<�_���mn~�
"��&S�fd�@��@�A l���K3+0�Ђˋ[Qr��:r���ڰ)���e�];�2qF\���劽\l6�ύ��X�<�CјhY񆕣%���a_����I�܆5G ���ذ0���{�@D��G�q"�(~��`�Q���|'1�T2Kz��hYp���@�d�����ʙ�� ����{�AʦɎ�B����1&%��|��D ��r���Ȟ>���5ɉ���7[����ᢹ�cv\��+�U��?��2Q��/z��iP��	𗩕��ꩉ����Joo7����~Ǆ���[���b� Bs����^M��ۿ�����O�y���ǒ	)�7��$�1�F=�+((����ƖF3z�S�r��@!������
+�[�G/����Zt�`�ҫ�~����{��XN�޹��]�jK
�U '{�]5¬�`��:�hvG)�3+b`ō���v��DD��`_���=�s�
+��D��%��`�~���C�G��?���0��G�5Y��W���	}���|�y�b����>��
����G��v�@D�.`����Ұ��Wa�?1�D�
�#P8��P���#���|����G�UZ�eO^�M����� }�%d���w�~8��#2�9Ye��tA�ukKoE$�6OZ�k�<��������D�#S�_V��PpS��i�ߜ?���D��:�ʈ�������I{�DW���l���M�1�	�
+�,�,��ܼ'�.���^N?����W�WW�������$G!"uq���N���|���x$�M�~�_v���ҳ�d�$-��m��=�#�B�_�[W�	E�l��!J�{)�S�p�a߹s�J�Iì�v�Z�����[o�e��^�S������P�jȥ!-A�P�D=�/[V+�� K��ג�g�S�~rڰ�ЋGA��1�r�$�����};P��j���rɹ��J�P\�2�� ��qU�ͽLb�S���J���z�;�������E��H���`��Q�L6& $��HZ���9?H�V39H+���0y�=���T ��,[����|�DD/��hL u�3@� &���aI�b[{H-�Q/�2>��8�]����?����4To\��>�|�U$}�N���R�=��G~��gy���$[�w;��8��N�OgN�J/���w{��kox���8! >�����8����0iϘ�\PP�xq����l����0A�k�R�5�H����|�4�mn�'�t}���y>ʷ��O�w���t������yk{ۍ9Vi)ƮrV��y�K��n�DB���smH�HG�>;�2	Y���
�枼T�e�E�!�wϐ��@� ���9�ɋ��9� ���Xs�)&y�\�)H��-�P������)2V�p��z�U&�����j�@U�U��q��Mf�6�A*����G���o�j/�B" �l<<�|���[�	�
J�<���� ���鸙�D�!��3�<��U8�&����?!�򝑯��I���t���ؿB����*��Pu��0�l�z�Z��z�|>B�3GHe�G�!_�L�e�E��7�6���:©�S�O��"$ǎ��O\J������_xI��!R�[Z���(D����㓉�^ֱ3A/�I�/96;�|r��W	Y�}2�'��j�h|Q�9�3��	�+B�/����NZ_���޹��ܹ�I�W?���{���~��'�2Y��s?+$H����m��s§䚳R���si΋� C[=}�"�J��G�o珫�C)BDP<�C�!9!"D"��_:t��#C��(PH Γ���Ř���F�ɊT��\�Ҟ�cLD���2B�0����W��P�X^�;I}/?��9�Z��m2�T��L���aŏ�4�%~t2��V&����|�tʓ9yt$љ?���D����s�Ͱ�)�O+����(�&"�S�!���lADj3"�#b7��{�.���==�c�-���"H	��TW!�X� �[{���g.?�t�������O_�җ��/��9�-q;aH�_UZ�?�����ǏBD~d%��P���4&��E��߇�w��ɇ �lH��ѯWJ!�����!y����V���K[�����[��������x�|v�}������4Nv���ް�(b+6+x�J
���_(��i��G�N����I�5��G-\AD�����B�{�ࡄ
|�?���'���� �|A��WP�a�9�0Q�گ�y�f\�ED���d0/��t�ܑ�VS�N�Q<�Os�7h���ɼz�'Í9G��H�bɷ��|3�������xN�����{�\;�*d"½��y�y��LDfDN[���L�8�OAІ����6m�bIS>���S����s��	���즍�m[�N�K� ��	���{�t�����/�7���t��*��Oz�RbE�'p."RP��Q�������|��aF�>�M5��o��8���Y"�YɃ��H
�=U9�Q��0���}/������m�?L7o�J�o����6�8=!�{�u>=T��dCy�Il&��X	�T�5�� 5(�ŅE�A�)AQ��0�8%݌H�ӌ�g�r���J�崣����GʅPH����P��G�˼}�u��b^��>V�`BDÞMDvՃ�r2PB����y4E ��;�V�?�qA���}�F�*�����&�ҵ�>�eU�]韇{T���e��,��>$�?�I�k���i'�\s�6~7EDH��BDD���I.��ah��*�ÿ�|������&L���|�����Ҋ�/g�b�vb-]�p1���k�'�J��Kiiq1�XuS�z5O�1�HKAA��D!"?��dλiq]��#{g�_��Z����RO¬�n�*�0�����u����V`��m-a�&K��]��������?�I��x����i���v����5�#�R��`s066Ca␸Qvl��bA���������AeK)�+M��l݀�d��'~��g�2L�K���`A���6��M <��ή�S��;A���������d�� �>��A�9�@��Ӕr��X9,VE�����>i6%��F�H�a��U�?���%̖A�L���0� x�?$��Uy�t���*�d5�~L����&b�H~z�0����ʿ�N��:���%b2�h41��K.u�/w�"cr���d�1+�t������O���/�/��JZ]X2q��gH2%}"sAA�O�r�j4:����H����7ݨ��5AV��Ø���}k]�q?
��;o����V �00��Ӡ��jK�q��>�a,��K)tCy����{(�aO�����vw�ҷ�����;o��7o�>xߛ�=x���6w���N��z��J"4��R�"V$z��E�!=�vkV���j"*J(�ss�V�l^�������8�'�����IT����A& B���>V��3�%�Se���i���9��!��'���i�?�q`(�LH�5�e���@�$o�.����,I��*L^`��Q�2Vy�:Q:����`������ڻ�*:�s��O��.�x2��ё-���u�����Iv�jK��AD��Fy�s�P��� �w���x�ɊK�-C5��!��tm=c�V�K��iye5�X>��y�rz��7Ӆs��ܬI_KaP��o���('ѯfAA����ς�������Ӹ��D���T������1�<�V����.a?��az�� mn>Lw��Qy;�����
�=R���{R$(��H
;oz��d9omfV�hֽ\HE�9g��U&L��U%��g��O|j^*�0f�
22HA�Rf�~��_�*�O��oW{�C��&2V�& :[�r�-ō[�����G�{�R~�)o��w���E�c�L�J�
CQ���T�/��@VOfC�؏pPؾ�P�rm��xP���k�K|1LW���Ye�
��6dUXR�,��~-�Eľ���H~f2#y�\���V+f�Hy�3d
��"2�ory��F�"����@,�,9 ���vj�.���/�P.>q�;�>�ē����1>|	9�� �G��4�_䋇�(gق�����|����>I!��a��.$֋n�ce�b���~�a�������~�����n޼�=Qx��[����*#��j�n�o�D��JX� � ,��l���Y)*�
V�����7�z������<�p9�F4XDo_Ϫ�vl�E
���dU�$+`�����L�џ�GN���gc.�)�i""�����J��z�-�W����q�V�������墜Sy N׊"��&��KZP��}��g�"?GrO4�Hs`��*�*����V�LD���OX�y��s4�/��K�'�(xg�kk<c� |A2�����2^ȑ-;_�ߤt���w9�f���H��C�l-����.������W�3O?�xؓ���L�b��YFX�#��ɓ������|Fd���-��Ǘ�c��$D�>�\�%��!�����������]v�e�6v���v������)?|���r`�h��&J����H���a�� ���� �tkG�+��Ƃd�>X՘��lu�F����T��g���1'=v��B%��0�����^GD��҄��׭�l=�Y(�{�I��j!0���uu/����ptO��������c**��arSɐp��`�H��̐o�f<���%>6$���ɏ�y���E9&Ay�|�HgO�!�1W�����P┌���Y`�ǵ®�sA��u�Snr��o'��p� y�.�=?�"��f~a)�?s.����O�3'O��ǎ��/�	���J��Ƃ����|zL�	r�\��1��0�Nc�Y?@�Ya8���76�5v��L���7���z�-�0�vgg�C:�H�j�����X[�1�
�ْ,��AyaQ`b��T����:CA|՘������_���+��B	3q�V[��'C��ǫ4���
��{5��Ø7��WO��"Nss�:�fgJ�	�+f�=	?(���m��g�	� "�xL^���a+�Ky2�|����y�"2t�;�-aq�0 �AX(>��w�e~�它r��_���@�*9�@��
��71d5�� �*REy�*�#�=� �1Wj��!��=ubM�d)-�Υ�gϥ+W��+�^IO<qɄ��2d����|���2/((��(D���q�r�Uƫ*��XLD��T;�BC鰱��kz�y�5z��@�����勵���w�}7ݿ?�_���F�v���ѾHIGD�� �-Y�
?�0��k���J�X�}v�l��/(�X��|�"�Ĝ��Yi�<B�J'��}Va�['��qL�\|ˇ�2E�YQꌵ�a�V;v��W�EF�,V�{L؍a*�R�|�j�n��Ed�R2�%��|!�Bd���eD���5ڏ}Y r���Ed"<��c�G,�V�T,�%]&$��I}�8LD�,E�aM��~8l����X.��URU3��{r;�^1�M2�c-a2��"w��J��^/-/�^4҉ǽ��'�L/?�b:s|���v���G�"Yւ�/"
)��B��0d��}~��G�ǹ7M����{�U�;}e�{�+% �(=�����F�{�j�![?=x��$�����Ν��0����������'�-C(]�6C�1W�3��a�0LQ�K��'��1�2�B�2�b��T��r�-�����5�>��z�EH�o;u��JtXd�>�k���Pv�
āUa�֪E>J)f�C#k�/ ��)���3��4�P����X.�?V�̫X�Dq�b&��7[=��`��Cz � ?�KD�?b��1��n���!�x���G��NωF��H�#�1�٤Ud���)�����<&d^��O�\HgN�I/^�����OhȢ��/Xu�r�!� r��(<�~A����p���4B}SU� ����-��W�)E��<PJ(�	0�߽u3�ٟ+}���N7n\9��=�=H���C�g����:����:�}7�K�2���G�H;�B\�a�+�5Zʹ�����7p��X9Pΐ�,8ۗ#c�׵%ʇ��0�2[=ڶ�0���[�E��T1�eL���%
�H^���/�J�!��+��b��&V��,> ��K@��V�������R�C~�)�}a!�R�p@<��	ͽaG�EP s�DDy� hV�G�O�TH0�� 3D�@I?V� ̸���k#ޮ�t;�iW�񡾕��������1��k'ӳ"#��z"���7�\˕�����˶U��teSA���|n��D$k�)L��O=�����C,�C��R10HaHѱQ���=)v��}떿�Ü���-��{?���*���K�ַ�tR��{��I&��x�GJRda�JW�L"��P)S�	n���;��x��b[$6J;�q�d�]k;���AX�&n��m�z�p����r(�����p	��Ѐ�e�7J�;X+b��{�r �\c+��I�"V�L����CD���H�cȆ9;L�յ�������J�)�TSD�	�	"��c&~r )�2B��+CG�B�����5�s�4ۚ�o��DR��"��U@�S�V-����Zz������^IΝK�K+
wB����#ߟF!"_d"R�a��~*�B�*7�[��pgD5��pS��M���K�(8.[\�ճ��z�{^�X���N����o�ٷҭ[7���׼�xks�!�ߚ�UO� �� t�tg�7$��a-hx#7H
�b2�6�ia�d&�ߒ����?��E)��9�Rc�퉒,�e8�V �[8*d"B����Uy�Mv��e���W��&�;���L�U5�B&"�+����Ī��M&��"I�B�p�$Uȓd�!m�H��{^i�L�"Csd�B8�Ѕx�>D��H [�%��w�,8!;d�
 �3RY� �*�&@��������O�=�ᰒk b;���7ÂX�<줲:v�X�p�l:�|������'�H�O�NK+˄lҊ���]��v��낂/
)���وHƴ��:V��.�<}O�6��7	�:�\5򱍼���n�"�qH�!c�H�ٺ ��[��;��N���u��nߺ�n�f��]+���-�!`.J��UX�17笠zA?�p��pM$�ә!
��=TP�=�A�e�'�JQ�.�Ǿ(z����G��2�^�����Oa剸���Ak A>d½����V�E"�J+n��b�EKʟ�(�la^D��q��&"=��ΦX��.AB���Ḍ��fx�֒>��EZ�y��
�2�o��%�JG��ߡ����ba�"bvj�L�n�����ȉҝ��#���bZ^X�\H�"&�ϟK����}JN�8�/�fU���@�2�ZqTP�EA!"�>;yD�K7�Q��`I�(c��w��C��<[AUG�s)���䠬�D>��������6����nZ_�vv����F�v����")xO���vc�j��Ί Ȁ�B��E�27C$l���h��0���U�v����laq�=�i"����Y�R~+�����֎��Qa�2�5&�D "�����@(��%�������=���oXUD�  .� �� c+v�P��@��N���&���g��D�-��?Y�9-a!;2{�G�ȇ��u�8�ψ|��!"ܐJ?���<�#�_]�.6L��.�^�$���|Ixni*?�&!�O�N�/_NW�y6]:w>;�b�
�""�ܟ�?��((���BD
~��q�C��à���Vz:�������S�-�-�O��N��������(�Oy�p��ݣر0o����W��O
�	LjeNKf�-)5ve��ɰ|����D��WcM�|�������� =㋶�d�w. !��|����2�LH1<���@HP�y�nm&V�jL�̒$q��K��[YD�MR�1w_�u�5\��$C�@a�E옫9Ê����� ���Ō��r��u����Aӄٛ���(<=',�ʇ��ώR�sk��;�*/(����ǌ������lZY]M�/\H�?��?���SO{EN��r�PjT�AGg����JF>�����4
)(�<1��$�5����,-���Jׯ_Mo���t��t����`}+mm�Xà�" (�Ņ������R�b��˲�RZ����xN�0&"�8�Ͷ�p?4��5�N��H@.y.�6<��dq#&�ID+z����c��1J�޶��삈�3�����N�"!���@D"" +f'T�yHE������c(B$�$+r "�Ȑ�^e?ј&"�l-��tH>ő-D�g�IBL���H��ƅ���v�D:~�D:w�lz��'ӥ˗ӥ�Ҋ'#��E����U��l�#���#�����f"RP�9�Q5������cn�+"ź��!���n���g�{�{+}�;�Mo��v�}�#,�e"�L��MP`��iy1��,X�(�Ɇc���֒r�5���Ҝ""^+��g�^+&"
cli��C�M5J��~�Ed��0g�2��8ag�^w�#DBD9  }��1*)��|�������CE"��sU*@6����d��5V�O""��r��"1d�{��$��U��OB!���m�gU�'/]L'���k/��^}�������jT�2u��D��lB��l=9�BD
~�Q�HA��
z֡&�Jy�������h(�{�����Y���J������ޮ7NK�Hљa��� Μ��	ů�X���^(i=�Dɛ����YL,0\�Z�k��tH,&)���V =�!�LDx"]
�K��G�҃�,[�$�A���v���:�?��J� !�ԗ�V� E��8>�H�\:������PVE8��p�<�g�DE�Y���0�ī����������@͌RW�$�)��2H��ݰ��3�]I�\y>]<uF�}�sO��9�]�%��Ȥ�Qd����v��s���6


~8���D/ua/-�&�G!��u��(W)�P���ZZZZ�����z��ݾs7����[(t���la��ڊ�U��`��`�(P�kK	��B��N~Q����>ݷ��%���x��{cKɑÊ%����jҒ���[��]�љ��Gq(����wH3a�d���,Ô��<<JI�f[��4+��a@q<�3e��G�?�<{��	�įؖ������nn��7���]�����什~7a��I�p!�?5@X�?r��������|�@��J�s�ZM)����A&,L(e���[��;6룈��J�{{{��3(ּ�(�%H���C&L4e�,�(~�E�Џ�B�;�V�D��M���s��zĜ
��.�$U��h!��l���j�0$?��kMD�q�/�!$I��H�������A~�K�q;��BA��M�'�������������6�3��~"	?��\��I�A��F�A���L���W�N��;o��P`V�٘?����9��a������eh���sĴ2�5��K���c��Wuۿ��鍊7n�7��f��������/��;w�����ȥ�|}��+{s
C�I���!�د"��Ӳ�bܛǚð�I��{�o(]�	�-�Xq	��C8=��`��{��&�͓es� �.� =ߥ�l{c3�5æ_�A���
W��f�+��A�)\�%/;��q"L�;�e���F���Ab3L������1(R4Մ�|����L=��'�!@�������Ҏ]BL������崲��Μ>�V�K�^y!�=!�:y:-4gC.����G�dUF?�(�����ȴ
�FV����딉������������_�zz��W���|��7�i�=��~��&��Rr���$��LJ���m���w +� |]w֊oq��5�A�VI@�v��� (���#�$����m��#�F�b����=(�JaFo�Q�:�ևH�!�����G�hm��� 8�Y��Mל'<9�������	�Af���`%��)��8�ꍴ����t�A��Kؐy5j��)���������K�o�L�~����[i�ჴ�p#�1���Vԏ SX��y���R<^"RP�9��9�� wR��G�TK~D�����y,�^�l���{�'>��$G�w����l-O����H�9̈�=c)5d˽�	P�!gV�V�V���R�&cr?�,�����lقbB#?��P(Y�2~bG��b#8#����qC�:f�L���d�"
�bU�ȇ��!��P�^�K�x��%��b���x���q>V��;�N�4���i�n��Q5tf�-�����݌�B���!>K���z�q�Vz���|\�~�_�f�i����'��q�!��/(x|(D���s�����E��h�u����}����owLJ];���_��nݺ��ݮ74ô��ǳi��LC�g�瘣�ee�R�� �;��DIe�d��E6�/X��u?<$eh���"�@p�����T�N,:�.ly?#��B '�
9�����:;�v�HH����i"ɊM��/��hz��>�*MUM�[�����7\��9�F&z�C�$"\~�-�|��>���싰�7�ݐF	A�ԁ�X&�+>]X&,>X��"��^'��|��޽��߸�>��Az�ݷ��$��To��AL��XD�;�ӓ]���?y"R�c��[պ��q|^�]?��}����b��a�{�h@~���n7��５n߾������X�lmm�>�scS����tRO��L��m�G�P�y"%
ͽ�i��!Kc+R��i��� �XG��ШHA��c����W��7֊��r�O��� (m�!l%�0�0�;�9��XY���&|��lT+H����?����o�px��#"��>�&�}�j0!Y�rDx $�����i�%���	r�`�j]q���|q���We�6�GYU�������M{�;i���tK����{����M��}�nz����Z�3,�|�ũ�

�qX�'/��أ������{hn�'��ad�[�r>6�I>��������*���~(��<?�*�iG�����w��Pa�vI�
�Q��aso�������}`Y��~ ����~��iey!��.�g.?�^~��t��zZ�/���%6>�[6��N��� �!4��.Kc¡>�ׇo뚿�U�49��_�S.u�\3SJ��!����{[T�r��_X ��1���l)<ѐԪ�[l-���*��w���س#���O ZM�� &��PS��!X��I�g�JvW�#��2-��[���ȋ3���L	�?� )�[�G���Ϗ�8��� Mi��pM]�	���U�"Ǡ6��2o�����uҎ��Ζ��t���t��5�����=���7����r`?a"�#"��ꢂ/��#���!����x>ʋ���y<��a��N=F��N=n������t��{@���?��N��3?�r4�ԅ���D3�)���S�3�} ��;Y~z��o\׹�vw6��g��/<��y�r:u�Tz����p���J'mony�*d����B��5;=p��?+E��`��������*ce�w��,�wQYWr�XD�{���-k<��o���;�����4�SS���������NP �����vED(+'��e"��uBBBv�r@�����s.����c��cc������}��"���ؽ�0�q��~�:��OÑť�o��3t�qP^�1�5ߋ|��	�W�B>��(J������������]��>�q�Cc�N�JǖWm}1����ǍBD~�y�ť]�95D�<B)�V�n|�C���ZI%���(Ld=x6��1��)�;�>Ӹ���l7���_�~9�gB��y�6�ALj����z �Qpx?B�	7gq�t�֭���o����ϞN���^���q���ŗ^I�����Ç���K|��_����V+���{�4�'�P)CǄ,��(�op��5D�#���4&=o�>��"K|���8)I��t��]�1]�{��x�z��(d2��Qepoݷ$k\�a3����Ǒ6����ȁ��#��*���u�3���ۓx%7�@��y�k�{T؇�e�:�9WXa��c�pEDt#>8(9MX*����En��Y����� wgϜMO��hy��+(���&�;�:����Z�i��W}������}��'� ��bd��~��p‴|�{�R��?��B]�y��� *��ѣ*�
N�~�������nY��x�ki�G���[����a��V�$l)�#�嘸�a�fuL���\�{��k׮�&�f+uu�|�ԙ����N;�~�~)����?x�$�_��2�,z�n���M��vj��`(I����ǺA�>�ib��EQ8�$X�˿W`�L^��재Jm��q��<�oLj����0��H��P`���4	���o�gc/�%�?�g+��=�Xg�	��z@:c�l���S�U]��ur��#��o�e ���ix&�Dy���76i�%I��í���Xi���_aRm @����A���W'�3ﱢj#���R�
����(����t������x�7��.(���V�~���	KV#0}�(���
�G<hX�:��x��|�A�t���p�9ܖ��g|\�7I������|X�r��c���������G���a�t&n����;|L���q��":~�TzᅗS��K7o�I�tܿ���}�]�^��z���g���_�������u�Fb��isk=m�l���wӃ�w�p�wgD0�P#�o8�`1慌:ؗ�M�8 Lle�R)��e�RX�m�7ʵ�@�⌃o���R9�[5AD���<�0B_�!��O9��]gϽ�*7�#�"[v����dj�L�����(��̦d� m
΋�OA��x�-ܧ,Av��Ga��ؙ��̷ȃ����d����O	� ��I�q3�My0�ae_>��m�
~b5�m�ǀ���4���>���?B�Y�U�cZ�Ao�Q�4�f��Í�#�Ga:�����8\3>*w� ;P
y������cn<��g����1u��K��:��QG}���y�q \�*lv�[)@�;*\�7a�����#C��(��:���������������Ν;i{k;�u��
�����rZ]^��c~FO
��<��m/f[p��)Iԥ�"�|��\��a�`�:I���p0�]S"A�pDs)8���wAt�7t�Xy��ʑ�����Q.�y΢��r(9���Qu�g�\�Ƈʈa.,�or��q����հTv
+��O��u�|��������� �J��3��W�.q�I�w�ܵ����*(xP~�V�8�x�~y@nP���������<Ý�4�>����r?���հyB�Ub^~G�[��N8~��$�ܣɲ�Ȳ#�H/+��e�ޠ��`����q��ǽܜ�K�.y�ݲ
���{��[�p��K�����M��W��/���,<�2y��CSC��?.�+�1�754���Nۧ�Q�H�� ;^�At�(��u�|6�+(��Hq+��z����!VN̤�zaK+���֦���S�����+�W�B��;�	���=rv�y���ڄ˪���Y�P[�O@0��+�U��W*$��W>W�XY�h�f��F�k/OU�ZH��u󧊊��������D���Η���-q�ЕO�y��w҇�����o�?��o������O�s�Τ�Ǐ�瞹���������?��ӥ'/���{/�w��t��]�9�pg��ٔ��������d���̨��!VӘ(o'uC���^��9����]���,�,�t�|�_���_���#��R9�M����e��!6m�Sހ�o�3��O��a�O_��gU��#���Ե�:�*9����	;c�;�R�.�u��`ĥk�XU=�[&[U\���f���u��#XN����~N�SaLʆ�L\1T� #��m�5D7ڵ�M�an�[h~Cy��~�\y6�Ư�zz�����:����?9�؉��/���\����LXiˁ_\��[��=�6��Í������/0ʅ	q(Y��D�d�B��|�2�~�lf� � !Y	�c��ȍDc�L��qE�BG����1������Oq�LYQ�g���6{�a�9��(y����&��q-�P�=+� 5��U��t����j���7^t��X���ߐL6P.A�5�&�\�-��iav޽�-��i�|y���	0ׁ��4ڳJK{6��@B��V�䯶���`j&o@���2EQح~ge\��L9��B���BE8��-�=;ħ��6�3j��G��|�;�AZ�+a ����Z�������� "1���s<���"%O�7��%�����gi��������7�Cyw�<Py+L��!&�[9��~l�N}c�4 m�{oM�[�5�Pe��Ag��V��<MDH}XY*"���f�G�������O��İ{k��Yڭy姼���dRB�{G�Z��Y��:"9Qd;T
�yꨅ���pU]g"Bf������_�N~�@�����B��dPܙ�d"Bx&"�3�s����(�	��N�����zly���^K���܇�γ8(���{��܅��+_�r����L:}�t��F�a�x�!"�@���fS��zlݴ����oK�%oN��L��v�������k�o��N,Y��?݀^�^D���O{���0y�y�iT�Py��M	���A��/��{Ζh�h�l2�}HAd/t��O^a���d�&���o�|GB�P>ȓ{��Fx���]�A��t��	M�"eu5А���=�d����Q_�+^��	�/��?�&��1@���Ѭ���^�N�_�A��(%�2A*�pU�|�ܙ��?pz��
Za揓��yCC�FS�<bks��{b`��9��!��U�x���Μ9�n߽岳��<�9M5��J�B�o�p�/�%|+E�����n�G�W�Ge��l	��7�zχ�� �	�k���H=�(W�r���?�ǿ�>x�N;�Ξ=��֎+m�ӯ�׬�����/�/'O�L��v��?����ﾕ�ܺoKd������*B��9%��j)9=d"7��H�+V��Y�ٖ�%Rm+�Q��i���+}̛`���ܜI�	+CN'ęg���Ԭ���Sσ !,�K����t)9!"���Է��Y��+��@\����J��-�\�A�d�O��<
���@�5����� =@¿����k�W�s?�k���$7�<��J9���""<�K�K++����"��Qs�ԙq�9�WA������&Q-s�xy2��A��WlW="v�d��+e9�b��8����j:q�x�CS(�^����>H�]��޿vզ�d�H� i��A~z^,s�2��l��˨�!B��#�^�n7�0@[=u�/[(�S*ܚ��@�hD䆗  !u�潲@����Q����Q4zțC�!"Mȱ��C4����R����,&:j�=�$��;�𖖖� ��(
��5���P��a':Ӭѣ�	$w�'d��U#O`��,��¥K����Ky�
����Dg@�܂��,H�ڊC^!�u�PGD����
&:2yA�kVzc�0�k�a���Ë́Ti���9���#C���p��z�I��z"ū�Y�Q���G���Q[g�;�~ ���?�<��}�+o�}8��������~��ߏ�/�_��_H�ϜH����?��/��b��������_���ҍ�����:�S�7L����;��m��E§�3A=9�,��Y��B�U<�Y�*&�*�v��9�]^��,�%���tU/���c�q��[�_,�����w5�DH�39�{<�w՝�����,.E��\ 2+�qn�Q���|�v�p���
���������6-G&���CU�U����tT/wFA$�w�S"���
�H������{�Nm��ډt\$������_J���BR�9�Gr���;m�>WA����\�����:����HD��z�ӵ�7�>�5P�2�U�duy%�9y�_�]�hl���_�u3ݹ/mn僧IPo�3�Y�� ��M �kF9�3AA!RӰ�hK~@W�(g���7���P	��1&M/�^?/j�����@=2V"0'�|��0�"�%=�7��yZ�E�,H�M��9!���J�ưE��aU�!c����v4>�U�&z,4N���O�qOA��&
�Ogbc+qz�$IM�� N��?�䑬�=إc+i�����;o+x*g�{Vʉ��Θ��hR(9$)�cDt
_e-�#p+�/���T-p���ϊ��u�hIQlô����*S���sҠT�`���������
�UO����d�>�J<�`�Y�o4f<g���7��tl�x��7�/I�IqP~gΜ�����H?��_M���󟦎�+����}��O�🦫�L7o�Mׯ^K���#�s����!ſ��y'����{���� c��Q:НҪ�ivG~c�\v~g�o������l3�H�V�ED��3�����C��[�#��2��r�8)s�#KCFژ\*@8���x�"�#���!d�=������S���Dy��i"B���g�Dɿ}���ꕉs:x��b�Ln��z3t�=
�謸��5?g�etJ����җ�������m(���|�8��ȰJ$*,��L5���*�9W��dPQ��a�K�@amlm���{7}�����~�}�خ�����N�����o��w���u�Nz���ׯ���~��?H���ή��=��z������v�;���IÎ^��0���t��A�c��#�W��� �"�,��4���L5(}���� ����������� �:;ݴ���?��ؚ1�5S&��/Yz=��wԋ�/�K���a�W���#�ݰ�X���FPDr�K�}�ۍ���p�����!��>�ɿz����1) h4���b�����\B������|�������
��Kfi9�6Pk�/�{��9����Ic��ٓg�G}����Ӽ=�cH�l����d���0�>���Q����[�q��Ph�u�<�
	hL��HY�c�	��aȖH�#�դR����S�wF��ũ��N���g+\Tu�2������g�} .���CJ��C��Y�r˅{�4�:�?������O�_L��\H��֟������~���姟J��?��z������y K�(����XXb�J�OX3���&V+�B.%�
LGWA�r_��mV��J�}LªVY�*��?�Q~x7�A�:�-��@TH$ǽqB湮��憞��q���}�j!��N��vO�;�:�a��� ���[�;-�Gʆ���#@z�gJ��"��M�����D�r��0�����J~�Ϸ  &�q�߸�h�������.'����~��.N-��vDF!��6ۭtb�	8�7���^
~d "4�4��0�:=^��u���G�OXa�2�,��^JOn��4��� �L��N����X����~���>H�o�H7�����,qw;��͍ݭ�������t����`k#m�yW
�#��'�ٽ5��VM���	�� �%E3ۯ�{{���zR)��f�2�!�������@�(L����i)\����!冂cR�~_9�F%es� �Q���+&��H�ix�D�I6��f�K�2P}m+Xe�|�T��Q*������x�@�J��8P� �H~ؽ��c��!ĺ�6���Y֔W})Y��d�R����#��n�@�U4�^����L~T��9$Lx�L=�||m-��K�R�(H�v^�f %H��ޓS�]_/��������������W#�5ʒ�0�4(r�T��K�/e�X��J]�hoGukWu�����D��Q9�T��8
����ʍ�J��|������$W�''�	k�Y�"��e�s.�ɦ�>1 �<�ɩ�=��J^�1�����.�Ng7���x����C��<sH:�m����a� �����K,U$0�Ja���\(�O�SGH'��>��o��	L��pDN���R�� kd�D������u8/)d@qS��2���^P~�	e��p[�C\M�u�7�:d>�)҉\������{�0�n����d~���:���@���$"N	e���������<��ix�7i��a1dÏ.HA����@Ω��8�	m��Ȅ���Lg��vݲ>g��ʅw��E�,�a/5�>�={&-..��M��w�_���.(�<�w�*���?P��&̄4ؐ�����K�"���z���6��+4RoԦB5�4v4�9�ѿ��A셰~/}x�*vV���������x~n.�4�d�Ń�l����*\��K�֍�z���ĜO�S;�ٟ�a ^�}��z�d��^6/�^ҺҼ+�DX��{��;j��z��I���#���Mz�,�$<p^xd���{!�hȼCi���Y]�X� �SW���m��+���$W�%�}[+��k������z���̑�'�>�"�u��q�B��B��G�2X~IZfڕr��ZTٌ.�͵��Cjr�J�oav����V��o�N;;["�j��V�a�}K������5�{���z�[1�CiD�);�{(~�\�r�<�)c$e�v�ipE�LtE�!4�'?W�ͺ�ȧ�I.yht��ܪyh��"�i�=�9���%|�#ǥ߹l�{D�;�pLSe8S��J;u��_K/��j�'�Oҍ�7����ډ5�'�����|%���t���،�|�K�Ku]���[�w?��h������g�׋K���5��t.H 󍜍��81�#7� Q���s�#����.hX�DމY�!�YY6J^P>}�ܺ��_�y�[�=���_���˯eP]R\6Gy����k97)p�9)�qh�s�������P3ib����m�$W�q'o �r�"����F�F�����k�>)`�_���%���͵���V�)�.̧�W�M���_IO]��ZJ����(w�.������"�_�w��*s4F�JQ���y1�1�!O�M��`w�vU�������R&�����(�N���bN���ȟ�;V��⭱YVa�+����5K=	S�č�ޅPB�pz��"$���$�sW�5�`�@Ρ�>���w44�u)y)�:��B�R�F���踆�`��W(M��&��M�j�]�� 7�g�A�Ԋ7��i�h�P��E#�[��hEpo��͊�x��2��5Z;�q��5q9N�Ԍ�|rD�]ң�����ò��T2�cS���*R�k���E/�fe���UnO?��'V~���o��#�&y֜�""_r���������=[��@�Ő%0�	�G^��K�xL��{ _K�J#XFʖ��h�h˄B
Қ�PJ�R,
�F�0�d��I���� �����Xn�?���@&�^�[vA0!�\~FD�gҿ���e�!�����ƻp����p/ݼu-�<y\iꧧ/?�67�^�E��^��n\�)"�IַUϣ���`�17�N���9&뉉���9�fi-��;@���������N	i�;�΅���?V�POx�Q��ɾ.���	�;asfu �(@���2@��EDW?���f�R��P��gD��Ȃ��|�d�g�.��R�("�� ,�D�S�*"B9~�������x#&a�����P���`�]��)� 7�>JDp�����:&~�U�!!L$Ο���\�t1�گ�zz�gӬ�]�%�Ag����t|804������t������5lw��{�i{{7v���J��ӭ۷������f%ƽ{�ҝ���pm�ݶ��:�~�{ޮ���=��.-.��W#��S���hD���̋��{�d��y����qcL�Fq�����e反�pK�]��-7���
C�g������s �2cz��K�J�ٽu��_~��&d���5�4�z���Ө3�����<e����77v�������Mq)){�>��M��U�^=CC����&���$�^����$^��lf\����Gڤ������W��_
�W�9�OӚ�K++��3��x4��1��u����!|�c��7�n�E�Q\����pp_�ty�#+����5q�O�GR���&���=r�����QyB�&2����Z���B�q�r�y��6���\�p&��s���Y\XJ/��J����J��ݡ�O]�����t��Zj�T�_I��ǩ��a�ڎȎ��
ee+���W� e�4J&+F��$i�Eժ���H�)�(7����A]Bnz�z���A}�lܓ�����XY�Iڊ;�.?�4�*��[�p=k@��{r���k��o=��#�_�W.�ޏc^��'���r��ڐݐ
�lDg�u����y&�����NϪ|u�:\�����t_���뭞@�uf�=��=i_������Ϧ.��ϊ��3�������TP�#�Wb�
��v'�o�����{+����}?���F�w�z␊��������lm���N���K��|�-�����-��7�c�=]��ѣ��"����8����$K5���7�j����U�z��+���1n��^��4jg��9���}@�����xE~z(�0}�v���.�����3w���W��� �n<7�����	�'��#&6҈q�Ja� ����fvOP(S�
��4GXx�P����]7�Ѹ�jM�Zu�]�YkI)*�~^&U��Sʋ}$��-��+�Ŷ�4V�N��'V8�Yj�-�G�v���yނ�B�`ff�֌��u�:"���?�f&��{'V��?�$Ǡ�8��奼�y<
K
ه�Ԕ_�iS:���+�Ur�� ˉ����0��� �,"�T�r�4�E����[6y��R'vwXB�)��A�kE��W䃬aѠ;ݽ����w�;�C0^C��Hc��V~�H� ���|Z^ZE]D�ϐ��C�~��,�A}S��"��	K2�� UB��ʭ��ә����Q�+���F�r�9��}����>���a���6]
��yL�+���^d��?|4 �I�}T׀6��an������;��H�����^+ �2����P�D���N�<!,D���������S���8�D�')ڮ��^����nuS��
ڑS�5��{NJ�U;{�uT��	�î��H�������eŇ;�j���ķ�N'�DJ�F���U4�m����s"L��S���������)�T�Ƈ�����Z��TM����ܗlu����Z�����ܦ���@�G�5l��z1N�[��$zsaE!~:�'��m�_L�S:�x���E���3fiR�Q���P:D����;��q���$�6lN��A�������B�"#s`l�Q:�1L��McN:�|���8l��9c��)�})#y���2S�Gh�|4k�dP���������E���W�ɟ���s�������Q ��&=�/Il�������V?�nOH��-��H;U~�tbc3:�ִXJ/;Zs�V:�kļ��ؚ�3���KV��M3�|R�y��g��b~H�R7X�㐒����~�\���� rq('%S0P�s�<�J��8���C�F��xEEⱄ1��deV)m=�Tzy��wW�,��?T^5�"Ez![�Ҿ��C9aQ��0̴C'B�qwGdH﷭�(m��1&�3�D��� ��b�cŒW\�4e$�|D� ƺ�3���f&~����S�+�&�1T�f�]��l������H��\��r$ovO��?����՝�!P,��ŏx!��Hʴ���� �qd� :_5�m�w�u�?���Ιx�������^:�b���S'�\��@���6���F���&0����'���	�u&�S�/���"�j��;l(:G���sEn!��7�zy)�K�T^5�( V�6�J�2�{w��[��P��Y��U�%�Sf�s��Q�\�Ѫ!c�H�Z�a@���&7L8Did31ʏyXB��I��#cȣ�^$l~�����v�B��z�%��W��X&�5XQ3�41�%gGN[6/��6�lJ��7d�d��}�Ao�}.jXS� `솼�Ԑ�Vp��%PI�� ���se �D�6�XF�%�i�Bp��#% � ��ce��M�qT�(b�e�*H�=ԥ���E�$Iq`�a�lM2�0��[���"��`(��+���CC�/���8c�fO�T\��?���?��R��Kwa+f��I����P���܅1u���zcE /�jE�U@�(L�K��q���9�'�㶖���N?fl��"����+/����|򏪁<�(���]e���ϓW-�K�#ߝ1�{���:o4��;Hy���_����?o
(8�
nvvAe΄n�М�Η2ƽ�	���xwMd��40��5��O��,f�������<Dv��e��J�ӈ�*yrdB������.Wȣj�~�\>����o�S�Ӈpy���U�Q:\���X������w�䥒P|�#����4~�#d� buL�Gy�������8�
�[��}���6�`�|��8���ʓuë������O���%�/�m M~7��	a�s����y���#&����h_�n_�=@��{RJ=);\���P��h4��j����ꠁ���=s6Yj�7��`e�.���x��2K��GR)"����:b�D��o�Q
�o�^x+���(�.un>b��iu��LcJ�H�6��u4D�9B@��3�I'���[�Q�L���R<>�(��͑ʹ �.��d�G��y�,Ȏ�8{�#��$Dxd�^LyP�#?�;��U�}�Wg�c:{{+�B��|�\qxk�*�f$J�ϐ����S�|cc=ݾu#=\��6�������]+YI&
+�q]�̃�}��u�]���*9�MΔ�G�D��Q�(T�:��VKK;|x #�ic�u˗��">��Ȇ5���Ue&_BB��'2�(���9���4� ��!�;�ٳ缩�r
+$���ق�A�r,���&�0ɿZ��M�Z�fYXHˋ��.¡̙��p۶ʐB��2�ܐ��CI!�R�g��s���m!�����t�&�,��rs�,������p9�5��U�W���!�*�1����e�-Ǐ1��g�;�gJ	�q@����ɻ~s���owp��n/�W~y�Hm�.t\�

~�8Pä�T�A���zK�����f�!��HŌ+�j��g���*�
�ĩ�g4ȼ<Y�f��QϋaƏ��J��64�:��YU��r�F��D��惄�O/#��j]x�!%^z��jdh8QF(	ݰBF>Vi�UTC��Dl.�/��� L��qb�(�	�����+j����1�B䎞�(+E��}#�/]C"|��ɱ:<�D=Q�亯V�+n��Xe��Ug�%��VZ!ms*'>8�V������p�l()v9e���<�b�;������d$7t(�h�U^|��@�r�ԣB��@=+)�})���Nz��~��|���UO{��"����v�4A�5T��=�*O8([ʍ��%_��W�\�qq�eE}4P�D���s��-Cl��C &��	��SW���o���g���^Q�.o��L�[��ɡN!n�	(��|�T�G�f[�u�Z�$�W�_z�e�R���o���l+��璝w�1�!�w�ջ�_+s�i��,��xr�������HiW� ��2a-с���iwo;u{{z�z�O��P�N������j��E_$�ð
s� 0�S���a��Y�a$&0Q����1l��:��3��y ����&�*I粑_��7$�Ag�����m+@�y�?,�a��Ǒ�|A$TƐ.��GX�t���=�y31|B�R��.�:`Mý7��-n�^q{�҇�>�9V_�w~?u���t����C>r��JB��ԟ�2܆�+e����ǈDD��
��H//3�	��2Y��4�L,�Vۤ�����t�F�_&)RK��R�R6(�<5&�IAxs��/K�������6��JzqiD0��+<���2�nk{C�M=�z���Hn$d��^��
��ƓFJg�Ln4j4$Ѩ���sL���F��on�4���V�9��B�q� p�rLc��W�MS�_�����~���1<I�HV	K7�]��e�|L�d�T7���B./��7H����"�$w���Bc��4�6ѓ�c�ʈ����2B ��(���'H��Ǟʞo�x�E�)h+]�K��{���B�i��fB28̥��g� �����=z�H~��Q�����0����]H��i��4���K�D,�pYU�w�&��]��+�9�i3Q�aP�$߄W�����b�D"��Zu~��B���\�&_Q�䷕.a�}\^YL��l}τX�bvT3IAK�G�ͭ���~��-��8aM���!����Ʉ��m����z�
��	�
�!��W�{~/U�������1❤\<$��M��c�,W�	
�Ä6_�/���K' �3�p0��ݩǮ}G;?U5:ݛN9��i��A�
R����01Qz�w�t`��h7�ٝ�
Ιϐ���O��:m�n��T-�{(V[��Y8����{�k���� *0;�-..yŋW�����@@�P��ۡ�D��;9P���L~��̆7`
��HѠj�yIi���͆=�0��H��H�$�F-��ӓ�2ѱ��d(6���Oϒ��T�=o��A��]1(����qс�bwoMW�o(/�z8e'�L>|p��'�ir�����8��ܻg��sg>DBc?���M����KI���&���)7V:l�Q����'���Cz�_@}2�R@�����\�g�5�#�f�a
��X,�!�׮�jȱ�yu����Ws`CYzC?=wݐ�Hs�5dϽ�i�q�y�!�pq�5�
�w�{V�?���:��,[����"eW�òڕ@�@*��"!����A{2��=E �,���޴;�׹�~_�d/vK�b��^��`ky�mnʽ�CL P(���͛׫㚿/�����x7}x��t���t�����0��.}�jr��蒑�d�:���(k�<LA{A@��� |T~p7wFޭ5w<�@�d�{.��m#�x��#�QW��d�.��a�8-G���#���ࣈ݁H����qd�I������_��4|8�������a�ǾN�R/�H'+L�EWpUB^H�ƙ7��(,�
7)�oxz74vT`����N&���X�Uo?���3h1@�����b��zޕ�T�f�1<A+�xjtEH�v0�y��Ը�L�wKik2�҄�{z�Q�qx�G�C/�/�d�t���4!��Ø��[(�*������_d�g�z���
���8�&Q"���c:��!���U�5=^�̈́���aHCi��$a�����+(�XF	1S��Qu���}��Ç(fGbH7�,0��)�C:)sܱ�'��=�])�;o�����H9$rqq.}�羞���e�|d&>�/"{������Q��/���Z�lq~^=���-s�<�׾8q�a���ǜ/�],4����S�|�W��UE�z@|�L�3ĜI�� IF~�L��<�t�|+�J�ӄ�L�����ina�Cn4g����ښ����W��B(B�?C�(o�}@���:��Y(�cNW����*cg{7�la���-�{�$���M[$[{���4��*&���l{RR,��tvLB�t�:R^���;l9��7��Ɔ���n{Xk	߽���6��lX�A�X��|!+9$41�U{�62����<���A��餐m��pH��3��]����������|ͯ|x��+�K���*k���0ĉ;:o��*�������k�#~:\�����g*o�U���ni�r`�m�	���JM�o�̙	�!U�O�6u��ic����%;~"=}����^�$rd�s����-(�Q��9Ɖ��=����I���z��XeV���)�;o֥+̲�ht06���:���pH��?�����=�aVJ��	K3������( ^b^6"70������( #/5J��}�57;�*%�[|t�iӋ�a���ת�Q�*d�!0�IC���#z���U#g��Lg,�P��}��hHIW4t*)=5<jg� 2���å��E � C�N���¡�h�� ��2�b�f���&��*�$ƈ{a��k��4��L�pU�ٍ.�r�8���b�v�ô~�����}�ת����yE����T+��|Vfa��زGn�~���v�DZZYP=S�+_�i�g�8$��<�R�сx&	���k� ��!��l�%�3L�U��r�=�Q�<�#m���-#5���"T3})�M���R�J&�G�t���tE�`ED�Uo$SM$�:�n���p��ð+�|�dS�h�P��􉈵����t�Թt��q[[���G(;�{��/���3�λ��\��|6�ծ�%vӥY��r}j�	���S8H����/����!8Qy�܄%6�;S�U�}(۩�zF)�\��Unv��$H��W��x�(���#Z�rd����P�>f�}��G�P�Ս)؏���9\�=oT�=�	��o�-�҄�HcxB��C}��!�#����������#�&5L�U:��W���Q) Ͻ� �� #n�Ii4"([��%���p(z�&�JqK�=�B`���W�og�Y�_V�L���=&R�Ӡ����t|e5-KA͊��g=��8���^kX��uͰMS�{��(r�!�0AR��@A`���g�U�<��	}5�X��|�=+5M"���^x�
gV��V:[�r\�ݤ�"I�nm�P���u��u�
A* =y��G�I��ba�\��y��)�|*��F� �?>-��)_���(l]��DF5�����y�u%��j���W�ݿ��W�@d'>2��#�V�D������B1���;:(7�k{n�uə�Xz��a��͇��(蕣4�\6u� P��;X���U+X��Dz� t��a�++� #�C�O�Cӯ܌ޛa�v�V�o��w�\<��_�s� ��Q����>5��.��rp�yV(&���䭻]��x�!�1��$��o5js��z���������ܹs�ԩS� �1�����~��I��&�9���ԩYM�O�L/�OO?�Dz���t���t��Y�Ϟ��szO�¢�{��S������C�ʝg���/iew�0y���^��3y��ʠ�g��+b'�8�:<��7�.2=�;O~�yW3TNj�L,*��<�;��Fk�EX� �<��z��)���6�	����@D��1I5扰�]%ϴHě#-(����������g��JQ�Ca۲P��=nvЌm��M�  X���R�1J��0h@tА���/�����kR$�A�u����)^]��0��&J��_:�F�������x��J����[ÊäD�E�9c�OT#�R�������8�$�ia+�r� w���h*,�%%��xћ������x�Jc��I���fN��<$\� #nD�y�&��3�A�;��0���2�<�4Jְ�0�FqIn����.�U^���%�a,E4V�Җ��S�XJ�����245�t/i�&�I���a�7��R&q�jQ�0��Q>4�L���{|����4HÊ��ݻwth�	u�娒ȍq�u	2�	�:���W��5���{����ގ��-��dWL F2����@��C�ɶ�!)�*�qCYQF8�ޙ����P$������+������P����Zؑ��C��ޛKO^J++K�d'�7wӽ{���w����YF-�c��~��\�SY���*�f�]p����S�UZʪ�*$�����S K]�g�J/�� ��*7������W�U�!�,�����o�!1�M��]�]�С�
�h�'� ?��|����N�\ �@�rcEpU���aq�vD�&o��<���RWLg���t�9qr�wA�!�?8���t�LBx��*�뜿�*��S����t')�����!��� �iO�h�ĉ�/����o�����S�h$�P��6����((�Qq`�����GUpzqQ�m!��i��v����zm����4&Vnu�m�q�2TL�y��5�YP>z!/K�2Y��G�k�_��_r�q鬈P�̣�E�� �_|];�:����T'�|(1����\��OG���\
X�#C���g�<�^�,�~�/aӳz������W��V�{�C,����&hzy���`�x���	K�T*�+99 
Ս����G>�DE1,n�􇹖|�J��y�qyr��Ġ�{�P�7r�F�!��[\z�,;v��fyʹ�r[X�O�RL�"��˿�v�����{V&�	yt9�vɃ�Bv�������$a�*�g�%x^�r,.��/\����vʂ4�WG�%�R����v�ݿ�[���[��t��+��~�:��P���<�d�f�6I���@��C2�*I�w:(�x��!=�_�|G=�Y)605=���Ν����YO�=��Dx�q�q*��/Û_\P��h�Y�*��w���H:� G���kA@�w�`5����0��	�ǒH�'�R����K�N���,�zyy��Y}cK#K�U�&4
�y1�sm�%�;��8����ahO�dm7b:�z�q��I��9ށ��*o�C�R7�Y�wrܖ(�@]R���k�V8���qM����oI�<u9ȭ���%�M�Q��>u��z�Լ�a�܄a%h��q㸢~����EgB@������
^yH��p���W
�uR���k�~��<��y�rz���mE:� �l���(?���?�}7 �v��L<��=�WǕWR�*HD�(<���9P�q#�4��4� *5�xx�٣�N�G�t�E���m�o�������uғ=s�l��Y�7���1��I��Y#�J��0�����!���x۸��1Wҩ�0ɓ���:C/J��_���߇|�AoGa�q�@���$}>wτV)A���w� *55,g���{i����.fR埔#
�E�ё�༿�9�|��˪,�$����BIcv�b�7��(1lJ\�?����q����[�H��� ��O��@�\7�?,ԕ16Mr��:��wK����ݿ�r�O�.=�������Յ��c�,e�/�w�w%/
�9<;;[��ͩ��=jH�+��Í&H��غ�0�φ���A���^�/V|�O?����7�|�������>ݸqC�'ˇ%�G����[��Df���4�Uj�?J]a��)7���"��XZg��H$��'�E#�g �З�?��ݽ/�F���"ݛ&Ŕ)���+�۶+�P�l��O�=���L�[.?��J�ȴ��E��c�Ic�*9�vz�d�����/�y�Y*�;�����6 ������L�T&̣�Ya��DL� &�Wle�;��7a��m �W�I��qf#C�yٮ<pM��\?י��}���<�J3�;DE"-A@A��g�sx�3~!��5�""�G�`�3���~��d5[�"~ɦ��iKp#it[DY�V��eX�YG�����8t˲a��;���MJ���0�ADn
��}G��aA@Sm���I�g�kϋ�(b�o�����f�������i^ߟ_t�,��ȹ�3�F^�x�<��d8��$��w(�����^�Do�Ǝ/�fи��D<زZn ���0v;��C̦p������E"MN2C�Ea�ԕ~���nm*��2��I�I6)W)���y��*h�Q����a������%.��r�﫧8��kL�����ٞS�%w,�D��-��u%m�2K2�c�Sj ��>srϽ~��zъ���(?Q4��"f���9yꔭ���Iw&��`YJy��M��O�+�"t��y�a޹w7uD�v;�d[ZY\�7cΞ>�rz���ӵkwԸ*�R|�	w{k+ͱ�^���Z��+Ϥ��Ө�MW?�j���8�Jj�5߽w'-.,�ee��;��X�rѫ]R�\[�a*�T~�}���I��a�r>�g�� #��'N8��KQ�9u�s蹳R���^K�;��_���w�y?�߻�����?J�o�M�������~�V:��'�����ò�G�ݼ�n)����|e.n!>�n�J�ֽ�jcs�q�sG�Iy����v����ú��I�1�m�}��t��m���A�S]o�N}lω<K3�<y2=��S�0x�+�E6�cECS���w�Q�A�u{WyH���$ʙ����� �������uen!�`)O���������p�[�z�0r3\��<��ٓ��
�bU�C�:v;ź@{��C�|�w�����_w"�ٱRA�P��t�B^R<$��/�{�����4��h� A��s �~��.h�ȰeP�|�kϞ����'Y�6uh��֐�.r����Y����.�r������̻aUi����VM{�6�'=K��W���{A�U=_�L�uF Ru��򽩃��߼���{i~�Xz��o��o��u54)C3?. "�o���p˽UX?�"cLD��b?���+��$~��QD�#_g"��qf�z�4����~!#4 4��R%˩�kZ��LD<ac
&;��
?�&n�-AcB����ٳ'�}��3��SO>�N�8���XS/|�J�����w������/%�;JƮ�%�����H�}O��������s�����{�z�|�]k��_z�ʉ&�R��DD��{�͢V���<�l:{挕�{ｗ�޿�����Q=s�l���_J'��"���L��>|�5H�t����O���7!z���ӝ���^R�K��̚�ř-����(������aZ�R:yrMD2�O7��v#}�����+��E�gUr���������}��pႇn߾�t����������ܕ+n�|����|���tWʙ%�g�^*[u{����Kn�3��IO<�"u�	��˄i�!5������}���I����/��F���`� J���Э[7�	��gϦE�Ύ���;�u�M~�ҥt��e՗}+N����6˓��oǚ��b{6ݸy;��ݷ��7К�/}9���+�k�<,_W}����Cv7�M~�a���s�m�c��8/������_5=񹭺�2���?�W��C*kk���$��!�9��a��r`����\�z��jDbo�HBHE�A�Ν;cr ?y�!B�l�_ȆH����w������1IU�r;?������U�T�	�vF����B��H���V�{"��[.#���Օ��zH�� @�lxx_�yywHÂ�ZX�s���C^��3�6$��ڮ�&'�3源Ƙ.�s����Q� Z�ǊwUu�9:X���;�[z��.���[n�h���yE�`	!~�[N�T�Ж�ufvi�z�g%��Inde��:~jh4dΖ���VĄ!?��W����;�xya`G�����i{�Isk���s/�����*D��'��XDl̀�C��*�{���O^ �訳(�*(�"���z���OD���d̈��S�"�G�r�A_��׃xV�`���G��I�Rx�O/�!d�ɗ?��L�qta�%��GW�����W^W~��x��E�l{A
���K]��^ڑ�ؒ�7�Rχ�٦�ŀ5�K_�i5�m5��֬����փ�)2!d0��K9�0J7�$��2|U�s\d�^/�������ˢmeXZ����u>^��I��{R$��P�X�~�F���?Χrƚ�o��n���{�ҍ�$�1)Ηҹ3RpjI瞈
����v��	5اݓ|�w��{w�0X=�2#�����ww9�P:�7���~D �٥���lX���L)r��?�1����O���^������>'�u\2QW�����a}XP�<���.s�����M�U���2�k�*�<iܑ��:�"%���V*L��0�<w�w��^ɴ�|z(�O�<�f�m-$�VJzNݤ�\?�&�zGronIc�P|+ʯ)Y���ً�#%�#���J��g90��u򡣲#�H�{�8�<�=�=���m��,,�3�>1�V9bI�PQo������y�z4.V���4�Iv_%���b�oKJ��P���X�7���M�{�����3&X�xw?�T߹�w)�k�Eo��0�-r�BgB�������z�mr!����"7�\��G,7�U����7T���kk�a�}�'��3,ISA|��'�+�!�X.瘨NY.P6�.����a	�ڂ�S?�i[��%�����ft�����)�s��8Ϩ�*.%�2�-����Yu:�}�����D��b��+�
)�\�"C�h�&���\U�q���XxD��"�>�M��Brh�a���	��%�[	��%��&��-��j��аL�4:c"t&U�9.�%�z�)��h����qϔ�Pq6g%����zz���i��|z�qW����u�l`��Dl��اAa򲳗G�F�1�F:L�|����# �a[V/�]���$f�PzC�í��Ə�m�I+�d�|g�i�aDv6H
�aʔ�I#n<�N�����VQ���1f39���
�￠l{��z�V�X²q��=ɰ`90�!?<�N� ���&!����ô����Ye�㲿M�ŀ���� �|��'�ҧ���n�1A��s�J~�4BbH'�vR��|��^=�v�9H����u�M�M"/�J3~P��]z�/���z|6�*��CI�L��7��T�]�o��l��/�p����G�8�3��	���Jg51�nK�����Ƀ��+~��e��ݖ�ސ�����Lǔ�&wRDX���|nnQ�d[yB�#�C�^Z\X2AX_P��G�i5g=��|�,�DGy�b��D9��(I�Q��\0T�������	�B���y����r�p��(\�C�����676|^�9�s"y���&�zh�2���	�	�2>7������p�Az��9!"�p��XN!��'�Cެ���[����k7�{X���c"M5�q��;d����\>�l�G���Az�_:N��+��P�wn�t�b t|��ԙh�h3�?�p,��v��xj���s��������C�*_����w��m��Xa�rfC�]u�Zjs�{���E"�LL����D_���������?�O�"x/U<���J�O�mV�y�s=�����Ǚ��j@��TʅƔ�Ci(���H��L?R���D�q��Ī�p��LH��{BDx��� yAuI��5���4��  	lxu��g���w���ȱ����������W#ݿ�Ng���)x5|�Ka���P$��.-���jhPµN?� �S��Ξ�)+���� .�l+�h�ǌ����Y��þ�B�j��HD��D��*�H+˯� ,AM��D�_P���{u̿�$��ʍ*
�{����ޮ�L阕���V]@v�V>����u'�mw<_���=P��I/�F�91��� �M�Pz(g\iz���!�F٢��]�YAF���;l�՞S��2� ���`�
qͶ���Ki�J6>/�EOk���������jwW����9C&ʟ�u(�������jUK,V�
�<���-�ʙwS�tAC��*d�_����D��.�h��RZQ��e���zJa(|�e��n[q�d���
�D��[�o�l���(z�7�V{�&r��a�����a"/���q��C��g/����C��s�s���G� RnLTF	�X;!�{�V���Ä鶇]�#H�4��쨞���	Ēw�:㉵rD����P}#+&|T�=�%$�sIԾ�:}�m��C�w��'��z@�R�g�o<�*;�u��Vn���T=�R����	ke�0i`�a�D|�����g.��@�!"��wz�JН\;�.\��~��������tUe&�!��iKj[� ��8K��5�$�����ֺ��E��{���;��[�����mOV�"���L�.���%#��4~��S
��8HD���'U*+&ϸm� �P�A��8�ĊH5��kzv�G����h����L�j�X�����B	�^
�K�C�A��������1u���Q����i ���Ti�~ti�Z~�*l�(��>��c庺O=y:=q���]�����e��I����ѻ{�����o���S�)Ϥ ��ê�	�N#zފ��U�2AY��0�9��F�;�vO�GZb�KeD+�sRN4��lH�G���� 36�Ĝ��:�hь�j,ջ6�Q��5�*�ΰ���rZ<)V��$�-����ߖL읠�-�I ��[�t09eUg�Wl�ި�0 d�޳�Qa�R�A�ā"" nh\sN�!�v��0~����x2�W��J���Ǟ7�}�=s�{k|�1����k����@�"�u��TgpOd1tCy�>H���=K����<m}T�(&�V����xNz,�����?{�'Wql�ݝ<�9�U�YB�($D���p~��q�~��8���� ���"���fm�yggf�;�rz�����j�ܹ�o��S��ռO
��èj#��������>�(�e�ɢ���	�a
���,�̤S#w�|,{� ���薙�Bjh ����ށ^����jak�����-��:�"%Jg�'�~(5d�fN�l��^�`�j��d�Ъ8��c]�EN���P���Dy�
h��}l�K��,��j{��x�����O�o���Q�5��ɾT��[$k���G���\���Sx�zf�Ex��	k;;�LMw�7��S�F1�����eͨ5��������3���I��K��i0m	�T4+/� /ţ}k��5R��>�l�Z�.��e�o�ة���Ȓ#s��fbca�f���l2.Zu)���Js�V��9YX�3 �Pf��u����y"�ʸۭ��Y�����&�%���ϓ魛�"�[��FLH2�\WHF\B�2��(����>�1�d�P�,y���4�1���hP�z"���BD��x�3��B����S�)��[�5	��w�G�������Nr�j� l1�d!�8es�����~�/�ƤI��a������z��زq6��m�m��V9�����?̉�,Aj=kH����:��兟��H��#�̕�J{�?���[�$�5ݯvC��+[����c���D�f]���%d�=+�����L�n��BHѪYE��Hn"M�C|��(�iUz��4�F��A:�Z�C�H�M��iOS+���j�e����HA��LSV�C�Aj[�ۑ>֡��J���J��$���(=�|�MI�Im��ַ��BĤ��+я~�!��
 ���(���C�)��6�h�w1n��V�H�ֵDR�љ�%��vP�$d�D�|yo�|u� ��K��&*���)�Aj��e_��rA�'���`�u׷̧��_�
ZZ���׼�|�?Ĺ��ǥ_���A�Y�;w�W��
/���Ϛ��?��s_��+h��3�����v�,\� ,?g9�2�(`e�cb�6� Y�X�V���A� ��X�����5��L�)�E��9s�Y>���"�(Tb@>c)�^4nƾ=�l|hzm���B܃��n�,H���`�oc ��?��V%Ʋtվ"���j���q�X��� C����ߓJ�$�#	Z���o�>TBR�)c��a�O�D�=~4�'��Cu��Ӊp�{Y~D{���i����s�ݍ��Z�w�}�լ�ƇXі�Ζ�������x�kc�����P�mC�6�b:V�y..'���|L�lL� Y�R{)�����б��ǩ�y.���q|r';
����+Y�[c�dz�c���n���D �#A� M�O���@D.!���)U�mj�"&	[�+ "�-+� ���D�b�Z��(�,.6�a@� ����lX� UE��S0Q5�S�#!���������Tn6Ԕ(�d*�֗���{�$/bq?F�Qs�[qp_-륕/����aSKV<G���1&�(�	h�.�.MVV Y	l�1>:��>�e��ޡCmk�yX�l[MX_���#�E�8���ڄ����
�ba����+��4D�	}jz1?�����<oB���mŪ��ޫ��*�Z�b��-�O��Q#����Xlc�Zr�%�����F�:ġ1ߘO"�w�gJ��c�x ���rZ��ʧ63�R���^�4��\s�F+Lf!�J y��3=o��w2=/p�~I�(�f� �X�J1�ѻBD�(J0Y���v?ǆ�PI��E�S�W�TcIx��CB��3���m;0�ׇ�1H�[q�����?f.I���`ێ���+/X����W,Z�*JQu�FIߓ&N@msn��'q�Gn��g��������/=���cb[�T7�(���+�����^�%�D0�-����j��qWׄ����T	]�	:�z�H�֖�+oP��'j3�R�
�Hp��+[m�������&�Є�G#
sM��(xe=8��Sp����Tq<p,y��Z=�ҋ/����@�-%��7�<�Ѥ�������>��V,Ǻu�p�_#di�pӒq�)˝ľ���2+����5W�TSJ�򲵣���M`M:T{���m��Ι������;wn3����W����N�Z���G�Ǹ�>*�-�N���P�W�I�"5�q�56&���Yv����w,���Uv)�g�:<Z
��1��6>�c�����̪��}2�%�1@���t��IP8�L�df��v�y.şLEs.�	E���Cm/"�(a���m�B�0 �P ǆi8��!�(�P���NĜ�/�J�j	[��C�7	4���`%>�������6<d$r$�������A��"d�f�>	 9���яb��رc�-�Kp qI�lw�i
WYC��4QLb"�w���Qy�V2�b��LV��PA M8�R�㓬<J#�(B��ꤴ�O_J��E��k�=���]�l끟L�0/�&�@jV.���k�6�va�6<���efg�PX�)jY�|Zj��{��y�(���+��^|�k�j�2�����ڤ��Ր�EIj�D� �L�|�@.�!��n{Z��G��� 0	z:>��zV������e�9��QU����w$@��w���N���]W:��ޣ���*��<�44��@��ޡa̚� �����=�\v�~|��������m8��{���~���V���?�+��׼�]X��l���������F>T��S��M��I"��_��W������_
�y��*,�e�)�ljQ���VVN�@�I �S4��t]V.�O =Ѧ��b�NWv�xU
�cdXш���{PW[���{x��p��Ȳ��G����C!�g��u׾��[I�(�!±�=x�c�(�tv0��7����G��0ɐ|�4;������u�p�۱c����k���·�i�ש���V��!gVK^�ePI�'�eѥ��]W�-P�$�( ��@͛3�@��ؿ7�z�	*��������]>o��Q�mљ�F��Ӗrj�" K/��)�U���f�1��Zu���\�I�-@,�Y�K����{�S�l�����J<O��$�#L�:��+O�wb��5Lu<iy�c�ȭ�23Ohaえ1ޮi�d�|mh�} "S��D� T��>'���A���y��]��9D�$ �A��a�@"�
D�Lj?R�g|J�C���2h�Ҹ�TN�$��C��PT����,�t��<6��>�];*�}�^��ɛ_LJE!SKV�H`*���-�W;+#T���U��H��y��=�8�66��Ւ	�<rݮ�y�%������z��xɼ�^?�������?�	�<��H�6	��}x�?�k_�&������mXt�����;{���� �<�x�Fzۑ����3��]|�%x��ߏ������UU���>�O~�SX��def�\�x����ߍo������#}��Ye�e��'?�{����w�	P��ĲI' "�]-�)<��0~%�:���s�?J��<���y�)��y8>BqZ��sޒ��ĻU[5�oN�_L]�,��h^�!�!F0GZ�z�yO!��o��+�@sK�B�y�7������j4���w�Cݸ�����yn���b�o�?�1y@7~�=�ٻ_C���E�g������.��h�{O������b)���Zޛh�y�SRz�~C�S��T�ĩ��FV.�Gb�%=k@��R��r����V]<�T��Ҳ��ݻ�� ���xt�b�L�2	�Z��͛QVV��~�K�;����0q�D���c{��	����������=G�H!o������7�q���j�>T��.��MM*=�HS4l0���ϼE�c��:u�|Wd	�4�VDI�Q��b(-=dS�R괯�@_����(ʱ7}�T<���xb�c[�6�vU��*"K�����l���i7�Y���5��M�	 ��js���%XI�i��B��hy��\+��٢ ��Y�� �M/��JYG9�j�0H��"OR��Ɠ'Mµ׾��&g5��s2��ӿD,�*oQ�H@��=�݀5�؄YNY˱���夥�v	^BX�f�z�������0���u�\MC&��h�����z�6�7�:6`���|�O"
G-���.4O�hN��t��8�?HfHV��������M;������Đ�dEuv�d46V�QĺT!��CQ��Q��ޭ;�=6.);��d`B��_T�(٣<O,?��y��γ΍�\�dp|ovn ��<y*^z�쪭ÕW_� ���>�)���|�}�c���hhl�Y���ں������3���mw��QXR�U�g�j��1��޽9�Z>+���T��}�V|�ӟ$���5�	�PZZ����ӟ�v��A�������W���%у�*�a��p���_I������hx494���9?���H6^���z|R���q��w�S���+�^2A����D��2{�����!�5�˯����~�s\q����-�{nz7f͚���� �ły���3��n�*w��}����\ގ�5u&�1{د׿�=�ҝwpy��_݃�|�h'�Q�%\�P��*��6>���鄇Ƽ�l���'��ڝ�GҨ5Hս|L�m�2i� ����(z�"���M̙�P��:F#a�V��o}��v
����;����J\r����.@sc�w��߃�4j�)���u��y�{���5�\?��/p��U�W[��.� mm���e��>thIp�()�����l՛6c]5E��)��V i��|IT���v�{Ķ'������܏g�z�������d�)Z�WS��b���V�^��h[���5�,��Y�����?C��3���+��3�*?0h�E�@E>i������6���6����±$�P6�)"?����Z����3f�<N��Lo�t�^3=�	0�S1c�`vN�7��8q40M�P���&$%�/@�BLBw�h���C�"Y�'�q��!�a�Ait!:�Ae2S����d�W���\�u��B��.f��}����oU�xؠpEB��h��W����L���ҍ�_\�����w����S��}��"�BuJ�W�H�J$í�ȩL�)0&�<e�����j-�z�̪b9(?֕?�&���l���]�K�K�"�Ø93Vޖ�E�˫H������8�0�^sZ��p��?���{}�����UM�������k�?��X��|�;ly�v�=��jA��3�<�^v)�>�l,^��̰_�ڝ��w�7�XSS��Ԏ5�g�>����޳�^r	
�s���3qƙga޼���S3��h{aǹQ|[-|�>L�>69����]����X�W����H���]�ܢ�XG9WL��׭��3N^ʃ4����'�sr��A�_��!V}�yҖ<FE/���>**.CWO������K�!��{��9�ϱ�&`�Ip���w�C~ �/�s���yR��c�����`i�����kw}.��������w456ģpRp��$kjBPWY��6��td���NyY����뻬��bjZ�cO|Hߓ8�����p��E#�b���`>j5��G��_�_|<I��i8w��ط� v��C`�iK�@���J�m@IiRXG�k�*���֭[0�r�Sq�%�a�ĉ8Tu��J$���Z:�"W}#ˁ�F\պ��~�k_��h�g�O����LK��E
��u��Ӗ���4�V��Ndge����")�wK+���,0�)�D��(�P�4����7��Σ��r�� ���z&�m"[+5���|��ғ���]<[��PY04��6���&���)�_�K�\�4�Y^t�C�S��!\y���-2�$�<��CI�s2�����$��L��N����y5������s�3� &#&-����a?:DdGgJ�gz|ܑ�G���3�Q�-���3�c�L��� ��(�ʡ�-���OE^A���(�f%�{�U��~��7�hj.Xi1۴�J����|��XJ$���.��FT�x����D��~�S���=kSZ�`X��<�DR�	��{I}7>�����iӺ�H?BY�*�Of¾&��i��A�{�}���;�q<`���X�
�d�vYY9��ʫp��b򔩨<Tm���Ttvt�ӟ�,R�ұh�B�t�q����?�QcT������8+r�����C�.��~vN�Ij���R�l�z:�6N�8�2�(�/Ǜѯ����y�@6iQW�C��Pm������=�q�G?��������[����Ԇ_��<��T �QXXjQs/��
TL����~N��d�LFAy��#�!-3�7�wޅ��mp��8VF (xX6�H�M�8GԮ;�����StP��~4v��~�'�����d�iOjL�G�����6�v&�8k����I{rH��O��$��ӗ"���(U�Gum%z9y�q<����l��l}��nÂyK8���W*CCλ��e��9���p����qƲ�{��K�@C4o��O>��9��_L|����@]\\��K�!+3��sP�����,����Dsk���Fm����+O'�b��#����,+)6��6�9��n�w��/����ҹ������ޠ�TiG�~�2H� ��%�T��|D1P���k:�|��6V�9��Y=���y���t��� ������48dt-�+zO���Lo�t�Ed�S�[�K�����^�7�Ct���Q�#~Ȭg�����{ƴ]cN���ˋs�s� Y�O���Ϭ�$�x���_��]�ʉJ�~MI;���i9�!g /?�Y��z�ؾ}��Гh�o2�Yq0�}J@j^V�%�lG˒��BRG���0 A��03k�K�㵱�%��9Zp"�~�]�_ψA)Ȕ;�M�����,*�옚���Ig\RI%�ģ]�\�w��`Μ�Xx�i��ګp�u����߹�h��"���>�>�x��x�����;�u5Ud�d�0�sp�M7YT�j����:�4���~��ux��o��+���̙�m3�'֬�\���a<����:m:A�!lxc#��ك��.� KW�'k�Ǜ��✝���F:��ǝ��U�>>a:>��D������h�D;�	���ʞ� ��Q�nhn�)�NAQI>������@rc�̹x�ŗ���ݍ�C�!E�����-�q�'>���ҝ������#����������w�����_�֮~
���[Y�� �	˘���,��J��%����	�G�D��U�̪$���uQ6I��!��3>��E`W�@]z��m�kR�щ��Kf�4��]�́��g�*��.�n/��������2/z"~t�%��Wv#9T��`>/[�9���Ʀ�֖CCr�w|=���2��5��Pm�O:4-#!��|9�XV�yY��*l��;v�Ɖ�/ �l��Ƞ��=w�]�U,�����?�ʱ�U1�D�)S��\��2�|��̿Û_���]���`���1k&�Ϙ��Ӧ`�ɘ0y�}�C!���R��CVn6ҳ2����@(���t��Q���e�S�b�(��"_9�zx������Aj_�Hϴi��G�C-'�[#�j�S��	A��I����ǔ57�%�6GOz�4w�W8Z���=w��G�'lGI@�Iq����ݦ)!%���#�A���Vht�htS����Wjy\��&C�DF��BOa�S�go^ziښ{�PfSUZ�A��)%�=�M�*B�C"�Z��!�M�XxH+ؑ�5�b@kfrgA�5?����s.�G��b�2�R��7����㕗_�=������Vh̚���x4YJSf>�A�g�Ư~�sL�15=��Ȅ��z�)|�O�� ���n���K�q�n������-�-�[��0|�$d�����߇e˖@�Ú���;��N|�S��s�?�'V��_����%��X�pi&�	^y�1l޴�^�]�������X�z�E��TE#�vt(�I�#�(=��9w,aN߾��4FA �A��d���J�U�[-��8�c�9�	��?$h��r$�YI�����i\U�N�Mz6q(	��&���HOڻ���Ǥ)3PZR�_AGW�
���)O���Y
2����R�?p+�=x՚��^��w�t#���;��ލ��'��}�C��f����Qk�/�x���E0о%*ױuw���6�Xq~I�R���"�V7~��ߡr}j\�ӮI�w"��8��3�����g��
�'����~�����h��G ���ą���MS�� 䠴�!�@(���hl��Ge��BAa&N���6i��|Ɔ�q�ʕ��ڧ֘5����6�ܴa:Z����,\���(��@GG��Q!ߣ�{&S�/\�����_���+���oc����3��\^L�4/�}�v�0�.�گF�W��١j
�Ș��x� �uV���Ķ��?�S�S�s�\��οi0��shX�Xs�)��/'9��I�U��om�IB�����C3j���g�M������~:�"��ck��{���O�J��qBȈ��ؼct�X�.��h�"/�3�H�W>�f46�MØ0wQ�
F$�Nll A���GV���w�U�#���D[�+j�(�k��RFm�L~a�>ɼ��z���+hnn�����p�R،P9J��d�,{bp��*��HykKk\�˓H�G�h���oJV�ĩ#z���ZU2�9������E[V��̓b��E=����>�Ge����\�v4�v�߿�n���E󡈰�y�|����]o'�!37Y9&x�Բ/��Q�j>�X;�.�oZځ�M�y��W��؈k���i]�a,_~�1���N���a��Ũ��&�)�9�C��	�ֽ���f�Z� �JǴ/�t�z8���;��Ԍ�����?`MuH��
(A��r�U���W��+� NA�Ə�qe����\�7_��W�S��b��#&��7Ҡo� �������F�����lGlxcS#c������aس[7���^#�Tc֌i���$?۷lƏ~�#�U��:~�"p�����6%��b��@����D�r�v�':���96lo=c>1�s#�Dp��������BR ����
1�-Ƙ�I�I��Ť� �h	vWF�m_[�്xe}^^߆-{�eD9zQ���Rz��:��a~��3��@s��)��=vecԓ��a��7���.��b��|�C�Gqa�J@�KM��׼�}��ػ� �?h���H1�ԃ�oF���[����9y���DUU�mĸ�㥤�=}�طo�E�%q������˭�!�{D��6�o�F��ض����1&����uM�l�C�fI�8y�L�e�ڠ����o���l���K���ٿ�)^�
�|OzF6BAYMҐ��M�+�a��.Z	5�r��5ӛ���;ނ���Ł%�B�i�)��# Į���}N��t��^'(�:ڍ@�4K��NW�!@#�.ox91	�(/�C�Y�^#��I3F���q{1�ߛ�P�6����
dFt�Cm}}#�}v-�[�	\R�՝��z��Ye�v!C� V��S�����}�QU�u�Z�TF�����@�̯ιs�S}U���hgi~�z$F�Ds�׿�m�[�Z�px���1s��H�(k��{4�Fþ�h�ʞ<i:ֽ��ӣ�'KOͦ���ּ������~8����y契�ضu�F�Ί!���ŐeEڜ�7_��:�v�p�a�mۺ�v��s�=��^{MM-�|�`��
,��#�>����()*��y+%�s��
�>>
j�7�T��HG�O�#�m��Ԟ����%���Ѿ>y��e=x����;�G"�#i|�7:����v4%h]���D�}����v-^�x�/&ғ�	_A酅�~@M�h+>�=�"� UX�aҮ,=1j�#�'��������،/���ؾ�}���`����?4D@�q�vS	���vѧ��=�ɤ$7����F�y�xy� �- �(��_���)HN����i�·/k�ٳ�Sq:R� ���姡d�rM_���g o��ȝt&�'���I�#�`>�IF���z v4a��&�<4���>���,��x�0����+=a?��y%�p�dq�$gp\ �s�c����MРe��P�~�b���g<.9�F���y�g��N=m{�1& ��%p��;aSӧOCE�#-��ȏ��,ZL�^U���L�:��-Muرs���x�R������}#��Y{;
��f�#����8���VD��)n>?�n*J+0s�L*d)'
��|����SPΡ~g�,��@�|��ac��Ӷ8��N��X���p2�U�1S37}�c�i�2���. i�
,!o���5}�Ԇ{��{¹Hև12?yI��̑LL����',N"H�kT�Z�PU���a�w-�C�q����s��C!�J��?��`�K�;��;h�򵉚�9�S����kط��P���NX�8I�!�A�$9`��eՀ�A²�90�ȩG��=L������knG(�Ts��q�~f�f�^㛩�����<l�b�oP�ތ�{��;�Bݮ�H��ή�Ǵ��Ma�uY�҂�|�6��!�����4�6���[�/�Gf��� �jw�u������#��E�X�6�+.ǩK�����w��طס	��1����UW]�k�67�b͚5ط?��	�� 9ʄ�M����J�Mm���6˨���J�����Al�����p��E��L���sV�SNń	�S����w�o�X*�97�ȡR�g9�ǅ�kN��?:%ulR�)�\��u"�������N���	�C����(3��hM"N
��L�`K}��wڸ��c�᥵�#?/��S�v��`5��d��iE��#���K�4k'��h�e�5@�?i��S8��2D��7����~��� �ט�"�N���l�I �1/���@���Ϥ�'�>i�Ee'h�E�<@�����F8R(�Icx�Ib^N�|���q�Of5��o>-C'�Wi�cS�xw��}�|HA*�=z�:�M=�a���?�7-�~�V\}����{ߋ�7���n�6�,,.�駟��b��>l+�&O�l;�
�k�Z���q��������Q|�S��K/m���ג7�l+Ұ&[	%����	#L^����ѱ��C���+�9W^z%�+�;B_G���š���d��ӱ��O9�&  �3�r�Ǌ��
�+f���ڱ�q�
u+^q��M��%1_!_�=gO�fY��CHfz��[�K�<���M��|#Ѱ9U�$�PVV���?�����ט���6�6j��>�Z[:�^7�g�iPs�N����?��	��]N��^d>N��m;�7�/B�A�,�g%�ȫ|d<���6��.�7��2q33�)bd��k�\��^��At���^AW�a�
p������L�L
�$G=�B�xc��5d�a�4Wa߾-��څ�;� 8y���m�U3J-LLzX�o����؆�^}�>�(jj��}�ɇȖ��4�8"a֡�����ǖ-[Q]S���61
��oUW[*nm`�<�$0��m���զ��������I[*�ON��.��`F:.��J|����%_�iӧ��'�ǢS�X=^y�-��	_��ʦ%�G,}�K��hM巃����� �!P&�h��^�X޶�EU���3~�M��?�y�\�8N�ŗ_�O�3Hgl߶w���Xz�bj�1�\�q�rR3����gI�D�,!s�Xb=��XQO��Hr#���b��  ��IDAT�+�r1����;k.F�G ����s9�a�g�s8�>���yF���r�����E9�j���eX��EDl_�eoZ��8r��ʑB�M	P7� �����|�����T��H�� RH���[R�^��˓�*+��T�ed �K�@OZ�0@�^8)���(��'z�d/��������EGK���E{u��e15-==}<��")�ߡC��JFsC#.8������{vl�8-�-��-�P_��g�euR?�?�t�����T!�G�V����5�J�����*=5�&LČi3�n-���㿟L'�%G��'E���Q���M+�!��u.����й^7�ܮ�/2t��=��#�y��#"gY`�n���f1!�8�z4Y��ʣ�9���0���Xv���pS��:�ߵ�9�D-�5��y��P�RHjVŴN�O@��U@�����{�s	b5��˶�1�<��J2RS����5sk5牓&����'d�K�����)�|��UL$I�Z<��cނy8�����5��6l�=?�%|z��	�	�Y{�؉���嗖�(�2�Db<w ���[k$Y�Hd��tJ��8Ú ��Dm��k#+Y__?�zz��ڊ��.��y��,/��x`WZ3
�)|��F��������P�B��Vc�[;Ǔ�@�
v.Z�=���'>�t�HG�������t�.�y��fd▏|�~���Q�ڵ/�[���ؔٝwމ��>����д�T�H�P=x�nT�Џ|e��o�m D�n��Y��c�+9�H;���/�U b�2�� v�6���p!�^�����W�²��b���H�����f����v��0���eS;.��ۉ+�$Y"�t��f�p��C`Q���T��H[1�VIIG� $�M	�#�Hx��1Fp��9�X��z����ᡰO&��ј�q�pL���7ė�M�>��BpE ��� q�c�?���4� �������1�I֡�੍ �� �q�V�K��0���n���̋�x��X>+�sBضq
��q�E���k��=6��3<������b��������A�r\���g�q�Yt��؊�{w����Ϗa���x����ӊ=��tݸ��C��|5��"Q� &@ٿ� ��>�!�������!#-�&N´)��^�x2�L�kI��H��a ���C�ݜ����Š�0Q>�#��*ʞ�1Ec��t�mt�(���y��2��xJ�s�A�0n�jLx���t=�􌛜��IA6����B2�n4�7Qx ��]3_~e5���1�����IBͱ�$�i��?�Q�m� ���)#
t%���Lôi�q��RS<˖��SO;^|�}�5���K0w�\�gfش�^vb!�>!�!��ٹt�d���[��F�W[���n��r9V0�H|J�a���v��L�1�2�=:�Qm�]>M����I��&d� ���"ɚ�e^������7��}�y2;��R�}z;s�"э|JR�~����@����,RK�
�����v�&���hҳ$��)�n��_Kc�A)�u�ۭ���(>��;p���#x���.���k���1��C�M�E!.P�:%�7q$���k����� �>E�]��Mm���O����O���69�H �Dj�jL�����u	-���;:�O�\��(N�1�d�\����^]W�1�rh�7
r�Q��"�x9&N���|1�9��a8����ڴ0��h(�@Ƃi�x匚O������f�|A�Y�>�C{'�[i��X�!��9�<w�f`f�2G��ۂ@�^� wS�Zz��!ؗo��n/����hIF���̀�i��l��R*I{���Q��G��2��$�I >�)���3�-T�]��6��!'?�<�Z���%.&)~���n�'�>���<Ob_����sx(@��j��l?��h�@Y]�r�)S�H<46ԧ�%��w�(�rL
��^�f��K2�q��ơ��d:�����ǑDq䈒�u�xI�$��0&$l	�N¥ıCyHT�SBIK�$�l�$=���ԇ��H�(��!*O!s'1�c>�K���O��YhZ��|M577��M�ɲ&�޺m]��چ�Ȳjh�n�}*��;z8:9u�;4Z��=�@S�.PRZZ�`ɒ%���& �"��#�L(''�e�8���eW\�3�^���
�#�@zVQ��|��l��DY��,ĺ�2���������#O?�T���,D�OK4��J|�=�i1�.���<9HB�v8�����ڎ@���Ń�i_;x.����&Xa�)���x������Qa��U%m�����Ĝ2�������dLr��9���t�J�C�,�}����7��/��~���룏��rVn.�'T��c�BYA@A��euc[Y����~8�9ߕ�_!:HȨ��A���J�]z���BK���R8<HA�o+������܄��<��:!�<��k_P�Բ(L	C1(@p�
dN|���0.�x�b�����#'H�@R�O�A�`����������sw'�@c?����6ڊ��F��l���?��B��+g��^���_�������l|룳���3q�.8=�i��K�d5���.��"�L����G���I�U�S�̒ �&�3-��z����E%'����&;�AK� �0���5�?�1^z�9H-if���v���X`��z����9��bƬ<��������o�4����L�w����`��G���i U3�/ю�/���R!k�E�&�6�sx���rw�����t2��� ���2�S���1��|$8k�	�aXbV$gvT���
�+�-�mV����H�j�n�4d�F	鹿�!�rx8l/�9�R�ʅ�L���7X�#$���37����cd�j�<�BY�s.�!��E����[)4Y�$�Զ$ "Qg�C�O9�N�� ��a[�t�m�UV���_�����XPP���tr�cȱ�Z>9@Qa6
�1s�l,\�+Ͽ�����\�K�&�%�4QU��E�d��ȱ�ڻ0:Eqv!n{��q����;[&dQ�,$���ς[ٕTv�M����1��t8Ġ���P(�� �� R���,��-Z�@���|"J$��4��( ������Y{f�iX�6!t��l�DY���:%1UH���i�D��t-q$4A%�KZ�j$�na��'��^[&*�6JcHB0 ,X���u:z���m�L�:y
Q�E�Z�����}�o��W��( �г��L��fQ�e>/�(��ʦ�K��"� @�s�
&�}WJ�3���I�O��ʂ�6�{�%��PYi�T^������}ؼe��0ȹ���s�-�Hԍ��>j��։�T�FBF�r,\�`�iK��nw=~�+3�@^<�4D��H���ל��n �w�����	B�2�	�X2R�0yB.Y��[����|�|�s���Jp�|�:'SK\���Kޕ�`��l�t�T|��������>3?�J>qs*�Oo$���2�f��޽6e�����(�9�ݱ��(�d�'��vt�(�H�\!�����TĐC�H�� ������*^z�Q��0�ϐ�D����������v��:D�Չ��Z�ص�6����{Ҁ_fV22������R�1���G�U��wi\j<ǌ�Y>��P�fll�?�A*_���L'��V�Id��c���sc���d�[�2�g)�L�ω���X�O��!�Q�B���JH��囖���nfD1J-e���>o�6�N������'���,t��tj\�]�֒۱Q7��p�����i�Ň�{����MAC�����L�z���C�g�OG�i�HE�T@��.�ܢ���k�Nv|�� $H�e��6�JGVv����;�����ڎÇ��2�l�͞�Pj��τ ��64&��[�XG~�UU㮯߅�����w�87����x��B>�p=QR�:���Us�6��kt�ì������M��(l+�4��JL���J�(���\�����V3)��@GB�J�&@��@"�?O�#t�C�a&y�89B��$+�ޣ�̚�w�^��}[]��j�P[�/T�-9$�05QVo��*��{�#8j�j�w�~�����hجC���6g������媲���0{Y��IV5'��ǖo���+$�D�m�\�5���X{�����CS�e:�A�?##æ��k0k�,��Atu�;?�	���O�!��1����Mē�Բ�Q<�B$eMD;�`zR��!�8#���}�a/��S�����ɽpE:����s�.�{o,��Nǭ7���Ұ|V 3�c�p<hߙ0��
���1�9���>����>��0�(��Ӓp����w��׾��>�z��oF*���n��;E���ña�3GI���m�H�(ⱽ�\]�Zӥe��7:2�=;����|x����پ{f��1}�4,Z�����w�lUئM�,�N[{v�lݾ�]�8����b��䕐�f��K�ҔG�?5b	n�.�q��m!�Iq,o��9����$�j�hˡ���d��L�8��U�f�����_�wB���ض.�LT�F�ٳ���W�D�m�u�̚1�*��׳}�$�Êi@������!{�� ��VKմo����d�i�]��뷼���Y)8�1y�̝3=}=�#�l����ϼ���Vj�3���̩�p�r(:aҠ5�O�k+�-.X����/`���شu�� N��QVVB �Ä	6m#�}�`�}|̙;����38�p8Bf�f��57�4_L��v�4��"v"�1�L���8p��]C�jlķ~�C�ݾ�LQ�ؖ6��&�����k��9ԗG:1q݀������Y������d7Y���fx^x�����QQO�_eP~j��SBȎO/v|&x�8�ƙ?>%��~S)��Y�~-wOϩ��SY�D�6��`(�0W^~)�C���k.Ǣ�31i�d����A�>�/��8���n8�Ɨ3�qꚎ�8?����^r����Y���q�[������3Ng9�x��́����7l��G���<6my�}���{�m>21w�y�3����#XX�a	<����!$�����că�0ߩ>�;��
���;�Y0�ŧ��+ʰ��L�6ˏIYcIps�
h� ,jS Z�,P���̕ߥ,��>e��x�"�ݳ)�1����bޤl����o'��2�%�L��{�xf��(��� � :D:����� 9=Ѓ%s=�^����]X����Yy#-������g�m�UVUZ,�T�1!>( m<O���|V��&����_X�	'a��=0^���,�sYSǬy��Y#-Vk��i?߼?"5���1m�t�Z�u2�L�[�M@D�H)��J�w�"j��oQ P �\5/;�0qh~\��e��LD,�f�i	�~��д�~��p�C�MZ���y��Ŭ$|ր5F9�:���Zj�g�`�A���˼� ���V� �<m�	���n2�X�n#�M�B����l�1k`��pX��cY��������~����f��/,Baq	:(\�j��͕"#-��S&"7/Mf�����Z�U���d�,Ggg7�T��Z�U����@?�4�~�9��J0�pd4�K���KO��~�S�ݽ�v��;o�=��xc�x�nc��#��ȑ~�����S�E�k:�ߒ���@]k���e�Wۚ����d��Л��w��^�u8p {�춘 �.F) �|����1���h2+M<
���F.Z�a|R��ީ� Y����yy�
�F�2��P�&@�j*��9�M3�4�{s��qکK�p�,䦦!���U_���Rу"����+Z�!�1�¶�>t�$ �:;�;�����v�Q�w�'�G�N�k�l�;t��ZmeZ/���<U6�|��t[C �g��k��ʕ�t+{�Q�ݳ�٥���ㄠ��{gF����#��/��,�.�c���/������h*����|H�"ڛ��ft,L��GD؉`z�����qŊR�+�(�eq�! ��'�r��K$,Q�����14�b��M��S�����L��3w�_ą i</݅y�0ef>�;�P����Y�?<�nh36O�8�z��H��l�7o���Y2i!�����1����P�~�Q�Is.,����I��������:��
��G�dxhȂ��g���q]Ow��sp��e�Ne������4J�y ;��t�E��V~Z"�1���d�,�x�vf�S1���*�/��O���'Z�dz��c��>�Ƙ�GrL�"]3�^�Y�L��f�5��H������H��x���0�#;7��
�Dl�|�L�,.|��	>/�/�c�f��{��"�ʈ�ͧ���۾֚�P�T'j�dP�]�0�����]x�����b�'1��&1�������z����q���w����L����|N~>:���y�xX���C!��)>Z��G���n�)�>$�p��~j�g���_����J�<�
�F
�1
7i'jH�J;��,����u�J\w���|���,�9K:��+��G��+)k�c��ɛ�m]XI�x��l�,)_�wL����CK���o��Xy�-�3NW�?w4w��N�� Ce?Ms|R�<^���1i�D�q�(+-�i<M�iU������;*���@D�����k ��U�!D�腗te�'���)S����_���Wxxn?�������ʭ�%�k���D���G�ݎ?NT׿�����w(O)�~4���l$~Ι7�_r)�F�ӟ�J�].fj}�7�Cp� iM��d �-C��*[
w^�00��hb��p�p,E�$��46@�m�k���X���*���!䧏"�5�@R>ȭ���+�Ӆ��)���J�N����Y�/��F�p�jZ��Z�2�hr9�>,>e"�N��`gZ���J\c��� \�����FP&�)�$_3.�,r�h�?�5�אb|/AR����<��P�(J�V͈W4�4�g'Ǒ�k�������iin���Q]Ym�e�ʕ�qdwOB�/�J�x�Ȁ�,F��+��̒�ZS�lFNj�d�1�����'��J�����R;�O�࿟�9i|���r2���xNt�����æ`x�z"%�[B�r湝��Cϊ�����L^�W��#6��]ݽ�<g�v�I�L��L4HLD�(���4�����1�д�t#Y�;G���<۩-�f�������Ԣ�����ҸC&�9����0`��}���;������ځ���<@��\G�=�=�C>YYdb�d�����Ԍ��F��O�����F�!F���2�?�O&W%ς�i�&(�������t�1*����Ĭ3	BX����2��@!A��eU���ӭ�;��i8Lm��zFھ@_l��������M�Ǧ#��!G^���%�D'b�P��8�T��3�L�}�t��	�(O��X0;y/Y��,����z��ٸ�󑙑i���i��&Ɔ���^f�ޮ���8\S�ڪ���ߠ��I!={�֧-=g�uǁ���	�c�vG�S�#]�UB`���7'ݓ8�����Kz���������泥�hz���C��<R�Ҕ��m�����VƤ��n���)���̲s08��p�ewQX��c���5 KB��ZJ���@;�O���*pՅy�\D �ה�¡��!ݺ��?��ғ$R$\�KS�9}���kɣ,�R4x��FEJ���K�Z�]�P`x8H��\yv�e�=�O�;��X3�ư��!5%�Hw=m���7����yR;�����$������䗡Ȼ���J�~N4���/�7Y1e������"<4�v�o.�u�-�eg�J��'˟x����-Jc;F�H��9�[xhj*�m�6Rd��oQb3H�?>9N�ՈO��G���S'��;)�!�I�D��J�C�+b�����[Wtd�"������4T1<��2ࡹu9E�p {C	�]NY�y�^2*	Ci�d������Q�R��L!=#Dញ��|jMj�h��Ma!�LZ|d������EQq1�aj��E5kK��QbKe���^�Lۄ�	$	r}�P㡥�+��Ŗ�;��S�������kN�=V=Z=���M�AW[G�Ep---ä�Ӱx���ׇ��B����Mz)�%��N�ˋ�I�~h�0�I��գ����n��wO���L��Gp�N�GF7F���MK��(|�y�o�<�)��z�1?� +b[��r�)�͔MIs�*���9�U�9��q
l�V����+��VCy>Y�	�Š ?��6�rxۙ��r~�y}���ʯ|L�y�m��:���Q�7�[�SIL[����'�@-=3������W]}5���m�;��ニ OۧO�6g�w�'MD��eJ0��˖�Ů��/~�<�
Z��T*䊺ʲ�5����Gqޅ�f�D	F� �唲 jS��Vn���LKK;Rv	!�E�ՅG��H\ӑ�/Q���t� ���xP3>?g�{8cA��X��L�jQ=w'Fz5ń�����@�°'��RҊ�Y2]#����f�5���g�Y!��"�!�BJ��Eq��8u2P@���OA@��m��8#��$��d�C�n�BL���>H�� /���Iha�l��~�he�49Ȼ���!rC(�C�Nѕ�G��a�هɑ*J<��%��b?<��Pq�"3=H A`���l���n�5�wҔB��>*NZyEfƲ�"`���E�3��r�	��-������`Ƭf,�1)���jz���?�E��m���fz������GV&�g��`�M^
�1����LA*���:( ���'+�F�F��"<_�ϱn�������-2��|��UUaY'�U9_;S����!m2�Y��|t��-q8��_�I��z�dz��cC�?��D��
v#��N�5i��vG�� H��Җ�miJ�KaaAs���$�r��A9Q��8
²�H{"C�������e�r�d�(@�zI�d$l���ʒ2���ƘV/֡�mĈ_f�����9s�t���طo_\Cw�	?�Bu�?ĸ�G�����è��ǦMm>W�x3��Z���������"A�Wtvucp`�B!������W�a��x떭hj�fU���V\���$L>�Қݬ2)T��s�y�><�����+b^�c���	�z�͑A��&{=d�TN����
d� ��m6�՟|a|\��f�Vw�S
�RSɼ�L���̷d#�~k#����j�MΧ���P10�����F�	d���C(��4���nDc��]�"�fG`+�S���9�#D�~*�6&̙3gb���X�p>�q�u��*G��g�����E���i3��߿�:�6l F�⼋W!�@u]5J�'����m<�E�#3�g���E�b}���l�v�t�|�V�跴P�f���s���G@Z�"�dz�PX�8R��(�3��%�CG�*�7��E;�C��+��
�8�x��"� �J��$h�%�SI�̘���%�'�!�������s���$�I��ɲ`�#3{��µ��cΔ 2��P;w��C�a�8��-�h"T�T��N�y��twr
��F�B�'DS�*Za&��I��*�S����������_[6T��0�`w���Q�Ve�MNI��;����0�؇��f�yr:z�x�ZC1g��8�[����S����w��)VJ��~�Z~�r*9SH����$���I��Gi�Y�'�Y�%(���G>U@���ܜ�f�X���킛J�aM��m[�O�6�Tx����V0�2�r��-p!�:K^@�C<TK�eS#<��~0�?t�g����5ɱ���x2�K�5G9�������P�Ϻ���q4)13	i��|5�!�Xhp����FqI�Mkttt�l�PZZa<���ۄ����w�����>7���&L��W���9J���2cJ�h��";�
!�4>��"��9`�{�u�PY]�.>��E��p@�IdȚ3�梤m���4��!I���[�H�J	Ji�#��s(��\b��	(,*Fmm��M�Va���==��9\�tw�W_�����/�O���`�sx�E�d�Xfv�m.��|�B ����3�˟ލ�f���Ĳ��`��Y(y�壦T��j�:�zq����ޝ[L3��ӿ���zYt�������L��.b]�V�#��[�i�z����}dziF+�ѲT-]M$�ˇw���6��{����R���-Z1�`A4����gb���4�)�?i�$\u����5kV�������@��.�l:�Y��Ԗ���zn��#f�	|��L�2����W��<<�4|�λp�%����߸�[���K�b�r���O��ČɳHGMH�)�W��U��bB�YMCiC5��bo����7���ֿr�..,�ۮ��g̰=r^{��^T��?�v)�94L�7�?�o����R"����VB�iH
��~�6|�ӟF?����z6���uE�E�$��.����
|�#���e���x���a0)#ZEO�K�>�8��'u"-+�e�2��0�0in�d�Z�1*^�$�w����B�@�m���vޮ�ه���f)�3|(�A����:Ӗ�91�����H�|�:��|�<�j;F�����Qe�5�WF!F3���aE���?�[��8X��Ru�<��ł���D�$>�Q=�$��x�V�%�o�q�X�d1 ���A{k3b#C�8���{N��)�|���3����e����4�{{QW{ض�Hr%x�UI��?(��Ɨ��A�D*U�4[����j-�*BA)!�/+3����ޟH�kG+e9e_�����^�Nt�d����"�ԧ�Ss��F������	�.K��V|��q�xI�yQ]O'"�Uex�	S-�"�&b���6�D�.�C�;@�J��ߴ���z��@ �|U�~Y�*r��#���em��"�!#-�@���R����d��<��j
GM)[�5g����OL�t=ʁ$�|$�roJ�;�!X~Yj�KFbfFX�KJ�́L{5���ւCq jߕ��#�'A]]M�v����-�	�*M�M�@l�d
*���o}�O?����%�`c>��c��m6��կ�;���l�@�m�&!h+���։[?|+^[��B %nm���^��4�<�ࣆ�AЗ�����Rc �RHe=DCԒ���c�2�8����9kɅ	j�$|��_�����=���~�}�4�m���N`������'��lkM�9y�F���|���h�Dڽ�J�������.��BF�__��L���b�-8x�
�|�M��߿�l�s�e���t�����t3�����7@2�b�}WF�����Ƈ?�^[��8&�IK�z:D����}/�����SӼ��̛6m@[KN[v:���o�c����@1�M�;Q:1Cv���xR]��C�?��n�_��hnk&��w�1�����r�P2����`:��#/�5��30MG�4�ξN��}��"������>��X�(׬*�)S|����F<ES²���:&�k������>�1Ҽ9������@0?W�`J+��~�����͉?R��I����S)i�����������OB�u�5!��+.���,A��u��`ρ�;��)��
H;��!>G%�tmH*��AQ���-FA�×��e�S�g�N� ]m���j9��"R�<�s1�x��N�ܲ�*�@��x�# P$_'�B2�Cʝ�lŃ�B�rh�)2+ٔ�t�n,�MKzR1W�*�?�U����4���ɩS�a����4�.�]����&�f9�Lo�t����m�I�!c��� 544m��9Q1u=��K53���1s�P��Ft��А�rVMM��3�ĕʼBdj�Դ55�
�y�����������.	E#Z�5��µK@pp��C��X��C������3Ǆ�L}�Vb�}:�MP�tי��E��9������.�{����˗��ξ �a�9���J-ߜ��4��~�5�&�d=jjn2-����� 8����ǘ���1�\)������Ƨ?�	t�w��g^�K�m�S�>�-�6b����"�}�`�"j�<��x嵭رm/��lt�������v�/��PG<%k�'!//�̳�>y����`=�tt4�4ȣ� �����0y�t\�k�������5�J2r��u�4)MK����������Xn�X�H�4�9sga��y&mwc�����e�'ְ-����(�DV?4���PR{���c��m��O�y�wl��}{�g�^�ܽ�&��_���M@��(ǁ�퓄���<x�C��fl�`4�%�uʿ�8_��q5�}��5�u��á�J�5-?�3s�M�UW�����������ۊ��JXv�O���$�őױ�o^t1�-]�76���׬A?��	p�o~�����)�*��k��#/5"�*&f���;B�c0 ϐ�u�r�ԋ��L�>�k.-é����7���1�h7�m��&ޠ{�����-�M �(�I#?#�"�I '�s�-&��`�'�Y׎�.d߰"$�(�������4�1��+�� 
�Sp֜Tt7��O>�qO������k���7>E�?�w�Ǌ �G~V\R�Ҳs���%ޱx��� i����#h���C{[���J
)�{?��vY\�ꦯ�=<�dh�j9po_z{��ᑰ���r+p��Յ��S���>�h��.�@?��Ӄ�������[�}���-�hnh�OM�4�4����������*�T���?�L��(�YX��J'꣓��j:�Hp*�BO^��)�%8r(��x.��{t���Ԍ3),�{�F��g��+'=����fe��t{.��]�*�FNv��ǒ��eQI��l:�KMͰO�'@�-�+�	X�hhyh�Kf��%?����,Ӥ�D�!�ߑO�2c���ط�҄iX��bp�N$ 4�cW��I����5����4 ^�{���P�X웮��$�� �v�ն���^S��@Z�788d��+8�e_!�HI��7�%cѢ�d<+��+�Qx~k_Y������i��~����[)t�¯�+���<��SX������!y��'S;fŐ��`Af_�� �����Ph���Kqt�̱Cd`J����R닭[���P�ݧ:i�LBE�'0*�ǂ���c�.2�z���g�E�b�J�bvK��4���K��e�&��s�P�S�$%�>u]����}~~�1��Zlߵ��������z+.����@B��.��W7n�7��t���\ä/�d�"<l�47�`^v�Rj~�+�y�����Ouu5�{�y��|G��w��6m)_�w��F��z衇<%�U�GI�tH�8_��j���;F�B�y�T�M��hY���f}"쿷��:̛=�B�?���ض���l9�,���<X��^߈���Bmo� =3���C�'J BM<��-u�0��Gp�%8}��H2�)��H[��d�tJ�3�߰�GӸa���:<����JOE6��,*K��p�M�H:�-,��9�P�\�� �M��Q"�X
���uM'���g>���#��a,4�S��¼��P�x�༽���T=� ��
��)_v��u��V��q$k�,�oɃE���Ja�hlh4kĪs�5����mO��C	il�!/O�`��+Yue�S�i�U�F��e����������_�K�yʚ*�]��lY�#�����A�L�0ǵ,:�_{2E��|��������ܼ,\t�E6}���"��M$�'��魒�"�r���C~nAG�	���b2q�~�!@!���#�m�N9Y��S>��3���";/�g!�@~N>AK&��l�eed������x�s#9�|oa1�NBV>96�.�B�W�iA��2���l
����̂"�[�HB+=+e����! �ǁ�Ud�)6 m���*�K0�yc�D�
#g<[Ź81>%��y��-��M_�P���Rt��%\�4O���{b�%q(�ø��f�K�S�Nª�γ6��x	.��j�R+�����$cc4ڏ��JT�M���|o��Q;�B_O;Ncm�O6���;��Ky"�' �<uJ�K�0�n�)ֆ��O�4� �S90�7F��J�H�!wn�nϩ*6�Of���r��]]��M�_$��^�l���n��<��5ʑM�� ���>d[����=�3��@���V*�~��!�ۿ�M�l�>�˹�K���~,?��VSDا=d�	V�G���M�him���S����h�i���GiL˟ǒ�=�X���^y��V���PE���+0c�{�w���-U�U��ĉ��Sm)	KZ�br���|R��Ϧ:�t�m��F�Nl[�+��V�	x�2�S�i
p-�ʴe�V<��j�����͂�Ti�g?�%6lق�P��iI
!%��ށ���p¤��P9̛��S3Q#��=(�?��XJ��ŦB!ǣh����3�d�*Z�"�O����	������E�DF��� ���KEF^1�.8�� U���Y�?�t�7�%ku��{때'��"}�V�w������#�iI(��� ^y�1���F��|�ろ�&0�$�&��
�z�a��h!H0���e��L��cO~R���k�nxÜ��4H�P�"�������φm&��d����������9��-�A�h�?}ן��M���eJ�Ѷ���'_�5#S��hN+�H@>.Z-%@#��ʩ)���Q��l�'+���H���,@�)�[�N��T:�H�h>[��P �O�Ew��<��9�=� Z�5��,!vY8
0d��5-+�߄�n�V��%dI	�Q{�ʥ��A�N��a����O6]&����M�β����d��sp�L�"�r,-���l��2���������TI� 8ڧ���Z�����'�F���
Pdu����Q|3�ڜ�#X��[�ui�J��ؐ��BS4b$r�����6��f�$~u,�Y�&�y����j���>m�JK�J�p�l۲�woe�J�P��N12�Q�(D|x�u�n��.�8��S#%S��#�82�$F9a���($32�-f˄�̳^�)mlXTX�K.��d���<��VTWV��G�k�+a9)-)�6U�H���Ps꧆��w�)���S�L�{L��9��bwPr������)mq����9N�bx�Q=x\�5��!�T���K�<h^Z�'�F������fΔ)x�%��ƫ߆�g!= �\�4lܶ�V�\|���(5&K���6	��mx�/�ޝ�&ymp���4-���O`�O�O�L�*��!M:��h�"sf�M2�v3���ɤ��N:gy�$�XG�lH��M�F��fʶ#/P�k�I���iɳ�n�/⥗^�G?zV�\��)8Y��[w`�S�`ڬY���w�ɗ�!%=I�T�� 8�X���X?��aL����_U��1��o�8N�f82�>�GC�ATV�&��5˨�ʫ6�Ӻ9N�	0��րg�}��7H ����L�H!��QY��+��y��_�q�86��vב�q���Գh��"��D�w�(��ǛǏ��dtGZ���¡m/a噧"�JV{_'�� ��ĺJ��:Q hȒ�xl�)S&a��9��6�9c�Ѹ�r䖏��L���_F:�`��-����~8���3ǰ�&�ȳ��������p��6Yd�����Ee�򯸤�`x&N����r;/��QRZn{H�F�]��3�þ*!_*($�/�5��Yf���s�
e�"���w���{8�R@����g�w��3�T�X ��-y������K�8�*�C⫴o%}ס��8O"�/�9~1�8�t�n����A�2MV�K�f��ߝwKh����p?�����en��2QJim
�������AG�.����З����'�"�i1t
.�+QE��ɶ��/�v�e�tH3���9T�p��1B�N�9l�>��M�IQ�xYɀ�̢j�D;��� �~�=19��"%�»��n�r��	J����]{�ƓO#�u�ܪ��:6�o����Txd��Xp�2445�:����C1�d�Q�7G�(0,ZhSiY��
�$-i*��_N��Qj�����Y����f.�O�3
�*lݼ���i.řћ�P�=x�P�Q�y箲�E{�_����W^~�M���(*�1�u����۶m��={���a�%b�(_��:ɡ?猕c��EKo��f|�@��P(+�����#٦؜g����HL����~�>����G9�����
̥P��=C�Q�#>��[PSYIڤ�a�x	"E�*�,f�Y�O4��z��g�y��}M�h��V�X�O>�$���c�9�-"G���R�ƒ�/?oBA�ζv�ٵ�,�ׯ�>p�\�� � I�HۛZ1����~�Ͽ ���=��o~�u�^5�-_��G����'Dn|�{P1{>��5H��pr:�=��;F�ׁ��A\vY.<;%�Ad'�-:��h'�{��Chi�'���l:�����ѪIg�Z��2����:>u��l\+��c͓G-�MN^1�'��;����S)q�x0~�e���?��cpۜ�]a7>��7�����|�w�]?��p3O �I?���G���f����b۾�x�����S��}���6l�\�Rd��؟3w�M�|f�g�uX �����B�^�wSSc#���p��?@��S��ݬ!�����<Z�� tѶ�.�l;ܓ3�+�P
hIQ	�R
i*�Κ����NBƫ�2*>�l�;��v�L��z"7�	߯�/^'n��/q��p'h�aX�;�}��3g<(%��魙�a�:~<A$�������(��Oz.�l�YXJ��\B<�.��c��_���oIU~%y9(�/6�^VV�	����ĜY�1����31y�̚1S&M�Ĳ�� �״�bthM�������i0H3�����9VeI�]̦'XGg@�Y�ι���O�yM)8�L���s'�??6�� ����z�p�b��я���'�z۷�@*��1�{zt(F��HF��AQs�Uiz����;H&b���wi�H�M�Y�i�N� M�d�Q,��{v����ஏ��_�
��l c�5���p�;r��r@�|6a+�T��z���H;BMʏ��T$��ɔ G@��y��ګvQei�H�=�ݹ{����,l��Ѩ�D�\U|$��IX��h�i7��.j�U,爘(�BR�*��"#�� +��h��o܅����#�%`��C��9sX��
d��s�x��G���f�q�hI����9'�S��7ˣ�ĹY5���F`��g���f�� 9�~�L��I��+����q����<����o~��/��J�_fQ��1��b%���oS۾¦�$����r�o�Ϙn4bE��m"��Ս9�gZ$�tm�O��-#�K�a$yzQ11	�.IGn�0Ҽj.
-a��M��o~�?������E4=������ޤ��� �V�xh��Ѥ(�pD���_gL��eD���p���Im��./鞼 �K/�&��?:��K�?�֎a��!6�\y-r
�����[���+�ü�K�f9�R��9Fd�())�W\�3�X��#�N�RY��3f͜���|&T�###9�Y6N��k��͋�2�\"aS���a(<�:h7t��L^I�ä�>֧��ڐS;��ܩ���=.<Fy-f�V̐/��g�py��dr<e��A 5�����.Bfv1r�&��x
�K��|�lL�4S����Y������E��y&�Jf��N8��6�:�����&��J[s��$	A9:iR��F#��pZ��$^
�HV�AY$�tM�;A�Z|6r�򐓝o�23[�K!c�
�@&�	M�ت�0롥��x���i,h���O$1'�M&XS����-?�GA��6�l|���v-�ʉG���z�Ɔ��a�VY���.(0�������?��2���AR�%#s���PF��ܗ��)4?��[��AM3y�dg����v��p9�Y��mi�Z�<$gM9��,~j��ՠ9InMc�`��عk;�C/�d���p�V
,h�AZ����߿��Gm��jA^nR���Lμݝ���œO�AOo�iwb����`g�]��y�����m�V%����vK6�����Ѐ�n#�
���]�RY�'�o��o��~������,Y� w���q��7�>.2bҐ,g����C�SO=M�2�w	@�Om ��6�);
vGKu,��M�h���.k�R��k䠨���N:���:�!��^�`*���x����g��E�}�5oC�����e��ӟ��9Θ1�����E����@1O4ժ����&*Qw7iZcb�4�X���ls&ӔK2��0oF E�"i�
�X�:[p��.̝M�C�������?<�'�x/��v��i���v���:+iʢ����ߤg�S ���l6D�3R�4�ECE�3I��P}��]t)>~�����jII��x'z�h��#��������l����c�����^~�V�S�/V�x�A�BA�ӣ�K�,����c��ݙ�ev���R,]��y�B&����}"�JP�����F�����I���'���4|�N�$˯��E��v���(��'%��l,LPC�I@���:'ȳ#�P�>�%Y������� �����F A����%yhlpJ12��(�=N��r:��e����Z�?wȡR&u�9$�up����C�'�e�q��a�WYx��'����ISlk��L�$���Z�&��.m�YI��%y|�"djY���hX$G�.�GZ�L���,������~׹��T�ш=oQi	n|�
���!�@N�|b2QR:��|P�ֆ��3Ck2k&��EQ�-�W�c��j^g���pRK�j!���1�缙�pg�Û�
_F��
{����X�(R}���3�u�C��{�V�}�X�	�?�k�b>���ᦛލ)�'��Y��m��@Fmm8@^����� �	z���e;�5??�m.sl���F�`����ys���عc�	e�HhE֡��<��&Ŧ����S�^.J"�ƬW�����}U7Q�ĒB��hu3¾:�Љ������o��g���O=���|�_į��8�w�W?�|�����}�s�
���$���1�����������6�&�K�Oj��@���gN⇄��C�,��]w�e�7�|�M�TVVڪ-��ġ���gc~�V7�}��"fO8/�%��F_{�e��;_���z^yn-\�T�2�q���ڗ�fQ`E�[O@~F��̻{�l7e�O�K�+���6o�l�V���I@ύ�}�r��x��EQ�g,(D��$G�:�C|n��m�s��A�L�4}�]ش�<p��ӟ������)[�7�u���Y��@���d�䘘>}��*��]ş�T��Vn�SRy������em�M�捹0�3��U���ы��n�����G�K�����G6�Da���;�q���^w=>v�-8��3,�����!L)Q�xN�:�TTT���ܔ��C��5}&��I;ڄs2��@ZjIЃN��|�ҳ������,�2l�s���C�Vo��Xw5v� p,k%�u���aA�T�m��U$�B���k=8��S׏=���?�f����V�J��#~�d�&%8�%�ȑ�-��_��CgT�����e�����8����oq4%}�v~����A�Y�?�ØY<��K�)��m���gN�Z_�O-M�R��p���3n��"z����ےK�����`)�/��#m�]\PH��5�[ۣ�K �R120��aǲ�AK�Af���HԒIm۶��mS�0TO/�n�`��c�y�+w~w��g�ڷ��o|��x��?������UL�P���x����4n�N�)Gښ�:����c[���E-U�t�yh����oݲ�`��4�֖6�� �;�ŵ[[k�غ��e�s��4/��H v��*H-��	`��EPdG��:��s̗d����!@�7k��׶*�p�T�$���%�t��Yǻ��3P�$_���(�������/ �t^z�u�ر_���q���'z�z?��7q�M�a��	��95w�੧��ί���k�:H�K F��$N(L G?I��L:�v�{�9ێ��N����Oj&z9��������)M}&�°�ca�3-��/�cB�� Z����ýmطg�I����7h�d�D�<��>�w<Լ=|��Cwvu@+$d=��Ҫ�������6�k��H���}(�I��sj��$,XPD �E�'���@JCS��^�a5!��k�T/�ΝAzO2ٽ{�2oҒ�f�}��y9��{}#^xi֮}����7DMM+2�G�Q"2�ǉcy���'Jc��3>�q4F>0�F���Ɔ7=���e��c���&8%�kim�P�T����"�ON�z�|_�#Qdffێ�"NE��6m��jaAN=�T/�J*�h��ʕO�.��	�����p�����(����ׯ��I��vlx�l{g5`��C�,�[�ɦ��j����`��+I��k��d:��5J������9;��a@D����-Ա4:�88,�z��\� MȷDWK�j�'i��$` p��'��Ŷ�9#�J��Bȟ�tj/���H���J�!��Ff��A�^a
c�Qᘖ�Ů��c�cO����hjm���<OA)�QUW��}�ػo�1QEQ<���kp���+��e�]I-q�M=iA�I:Wl����P�|Ew����������C��?�K����f���؂��jkU������{l鮦d�л����v2H��X��O���_���B���SAmx���^Q
��PP&7�� H��L�Dr��txB0���%_�$�o� &��syC�3�띟�E��kt��fg��ʗ�t�,���N��GMZ򣱥;�U��y�����/~k��:�)\#�|�4O���iˑUSR��{/~��`͚5�(�U�����I�� �h8j$HN� ��R�(0�S"��i3���1� ��G-�1<��;w�/]}b��Z1�;��n���a�`�4�}�N�*K =�H��t$�ʃ�
�o����<@<���1cr�ݠ�
D��������܅��\�e�{�N�5֠���]�6� (p�b!	�����'��IEp`_�o���=�8x���� � 9=S�X�(�BxtL>'G��?J���T?�3�l
x$܇����(��vk���Pd��F_'r���r���M_G�"��_r����U{Ai[�~�yY���mm�i�&���&Ш#�z��N�S�W���!:���:�����K)JAV��9dd�Y��m
BI��q̏�"��GX��=�
!��(/'��_���I��������9	�c5bG���ifHv�z*>-!)�d^r��5�L&��:��k�I���E��O@��Ɖ��抡��|9�,Z��,]��ˑ!ˁnu5�3ڇ�H����:1�_w)���p�}�����R�q����T�Ca�/gϟ���N�o܂o��#Զ�c_e%v��M&Ȓ���?��!j�;	�p뭟�5W݄��<���|��R;LӔ�� ����'���v�Ք���I��>?��Vo������ ��s�����g-��a�{F�2*�����g{��c]�y֠.-�֪'���}�n��{}l����;~M��eϊW���-
���ԉ	�8�S�b2�t,g�_�he`S��~DR�����p͕�a��r�A�M���ރ�*��WN�����4qX[׀��w7��������˃h�F� M����x,���mV��?�4,�����f� ��@CC������%h^�5}��H�K-��Ɔ��0B>B@,�"i	����+�
f"�BO�@G�������g>u;���o�r�!<���x��t�9N��*�iW��c�*f)蠂����p#��9ˡe�n��1�f?��\$u�0��+rDժ���2d��ע���M�=T�����l˽W�:�|!4�U_��Dc�E��m&�wb�K�>H��Tc��M{�h����s��՜�����#��;_¡?B�˷��	����RI�ОJv�#![*����(����w>�p��%��A[C3�Ø-ŗ���QP����R*�'<4lQS����,���8����c���؏̣����
��l9}aa>
K
ٖ�"Y+9�#�9�� e�%����9�Y��o�D����҉�M��I�)G�V��m�%��d:��'�1qD$����2�1���>�:�	ʱ��AzZ�!!����Vb8&�6����-�$Ð��\���7�����71���g��AK�=��0��9������PQ��S+0m�L�2�x,Z�{��óϬ5�Z��8L��q�Xв���c\x��X�a3����X�d��#c����26FGʁ��`�����c۶xj͓ذn"dl��!֑u#��t��>Bj���-����%D�VH���M���/GzcS��u�Ȃ"-�����jYu���Fv��l2G�x�)����������rv��.�ysM�)�Vh3���nj����Jj+�D�I����wS@
Px�;4F!<q�\�r�)�ǡ��Yi���p�~��/<s�N�_&j	�}FA�Kt��߻�n���g�Fβ�$
g:Fo����䤬���Gi��%��v�T|�^s&������IX��ϣ sEŅ�=w6&N�����M��91d�kކ)��aެ�8��K0�|���3x��'m_#v�99^q�e�jk�K��}����Km���k�G[{��:u���^�]{v`t(�Ύ6�ut�%���X�T�x?r�8uQ*�ʀ?e���a�gh��-���(�[�w\Ϛ5s��C=�����`ڴ�x׻n&ͤ��B��4f��~�a��akmM��32��6�>��g�ZDz�í�)�	���C"�D��N2@�H@t��#<D$�fC9I"�w,4@$܏���(Z�����.T���R�~� �m�B�2�Q�Sm��*�K>[��2��,2_����iii%�G���/bϾ�k��oh²��"h��3�ET�X�"dd|d ���ߋy�����\�ke-�K	 �8Φ`҄)�7w!�ϞG�R�Je�%1j�Z�H�[[�L'�?�mo�$�#�f�L�٭��3�4-ʕ#Ifm9�ie����8-�4 2��A�R0(I@�"�e��Z��x)4�d ~̝S��O���'P����9S0mr)�=��/��,ss��I�*?i��I��p�b̙?�++�E�q��硲�Mm���X~�٬���V����]8x`���J��g?��q7���E-12lsȲ���ɚ#��������e����~,ZF*�_N0w�\�\���YhV��.�W鱩-M��iQV�7��8P�D�)K��T���f2�HD�&�v�#]��,�=�8�z�)TUV�r��\������MI�q��%I�Ԗn�S�X�k��3������)�R��֌Y3&�Kp�B�  �k?5O�D~a!r�}��P`k� �����x��>�	AYE������mE�+�W�phP�q�A�5��;�M2�O.���z���=����y��'�� $H}�=س}\c^�'W�D���5�y�/pǆ�B�C,�~|��簑�US!rjԮ��-O�EL>4�����MRP\�+���`<��`{woEO_�M_��󋖇0�܏T�<���0����Ͷ�He�!s���%Mp��g�'���Na���V��.�k<i(j�H����d��RS����D��zV�V��$�U�����).v� -h�N�:STܬ��p�������(Z��L(/Ŏ���ޟ�����G?����:�C��'���O��6R�E�8��T7A��P[�;��l�j��� 6l����� �	��UW`��X~�E8mٹX��l~�$m\��r���*��g�v�9�"���r\r�������͞��w�,�,�LML�L'��Lz�YDl����+ip+b��e�;�U�5ع{�b��g;�g�������IP&b4������3�̙�7�����LE%,AvN��!r��� �̙���.Ayi	j�j��A�l�,t�t`��8B�~��5U��8�y%�vW�/-'-.+�|
�m{�a��g�|b9���"��a��X���I�0FAE�m"7Dͬ�����Z�b���vn݊���d���%�V�3~���x��9�m��D
R�c�.�޽�<�,�}�y���zE>5��f��	tK��{l�O��\�җ���3�ګ�PWS�ޞ~����$-'�C�c��m�R�@5?M��y�f<���̍9
\�g�ߌ'���t/)�ٝ��e^��:,Y�����~��4\y���x�]N��h䨨ꉎ���G�]�M#����֝$�-�bG�VQ�a��0�%=��������]�%�P�^;VE������cvf&��������e�X״�T��_���ަ$� ��W�_[���_�k���Gĺ֢���	��R�vc�ܻ5�j�z��N�Ȫn��?��$_��J���LXN����3��]��Iaؕ��H:�c!D�{Q���gO@npAŽ`���fz� �m�1tut�+�(3G��_xٹyx�{ߏj���@f	c��e)jnnş�� �t��8�d=��J�p�e�i�L����ٟ�gNѺ:áS����G~�|� MO� ���g�ד�z�V�������'�6��� #'œ��Q�]_�بD�P�^Z��lc2*���QpFE?��ݯ=>[�VTX���rS�����޻� ꩈ��R�9�%�>c6�3�����t�q^�B�Y�i'T8xmT�JeK�ZA(�o�liU�@�+Y��Tw��S����RKI6�N��鿟j{&�#�*�O���%r<M�@�u���ӦJX�J�V~:�	S K���Bs�bGG������"jGL]��߄ISP1e,9���LZ�w�0w�hj�Bwoy/���O�(�Bu�Y���<��Ӹ�B��˱���8�g/Κ���j��)�v6V�|ED�6Uu��x�p�/���&j�~�.�g�wZ���ʠ��ЦqrT}��W�شi����m�f���-������d�b\R{�w������Y��،��`/���������_z	/����m����~
k׮ş��'���;�yO�"���`�UE�+	>i�d���C�w����c�Z����K��S'M�|T��Y�Q" �T]$�j��q�@5�v<*�!�{EjS��m��mg�Ϙ�@�>��J�F���Μݾ#Ko��JV�"�vA�������@$�;��j�G�RN�#��ug޲�47�a���a�k/�����0�R<4M�@x���uw��P�@�Ƅ6Y������$�e��?�)>���a��((�û�}n��mX�p6�[RCl#�E0�E�e�fU��㱭�@�~_�YP&M.�3�L�-u�X�p1�**$��FcV��`�lŇ�WV#���y������*�~ _��"���r,(@�����$)9�_2�â1�����ٛ��V(�6�7�g�Ve�������y�|�"\��3�]:m�(�p�`�`\K�����>�ڹۜ�_��xD]�Ӂ�!uF+�K�.[�x1i���CtD�&�X���������9��D�Q���t���'���?�޲@D{Rȿc㦍ػo�y�k��d�V��AU~b��@�����Ef\�Iw��s�f��!!�Cͽ��c���(�0�����vG�8T�����Whq?C��;����	��M�H��`�����=��Uu�R���f<d��7mƽ��Oص��U>1��PA�T�E��"'�Z�� ���m�&֗O��<'�~��6P�fY���D��m��M;�;��'D@EL�6���N��8��q�<�����EOےw4���8�G����´΢�VQ���ڵ�?���ؒ��Ӹ^aEd�Py ��Ԯ�(h�\�mH%p���p�̿����Y"���G����K�L_��ٵ-��B��0o��V6i��QU�"|�	���dK�c|ol#���QN�#�T�f�Q�{$�{ �����0�ɢ����N�fiG���1LteQ#���a�R},���TN�?�f�~$���Ƌ��qX�Ň���]Ե5�ؼq#�����z�j��>f�`�b^�����-�Ųx"؊w�$���|�����w:����l�d�܍�� ���*\x�6ݡ霤��c,I�E�>`��l9ZkT8ձ��h�j���%�m�Ds[�z4�֣������=�|����:�u��Fm$������-�A�!�[i��VĆ���I ?D�s�Ԅ\�@--����O��|���0��k}��I��Up3�\��_}��!�I��� --h
�x�SBT(9��O���=N���&�5�U9Ѝّy664�C'=�����%r��)����҃��F��	dc�|��tu.�A��E2$i���`OY��|O�9bji��y��������k�����d,]��H%8h����Q+xkK/z(��8��f�ftt�u��_�/~�sl~c�I7�>�4���6i@���'�p!+'�
d6�Gm���c�^}	��m��G���4?�g��U�I�X���
ɶ`m���BP��4j;b�N�u��<��m"	𙯃>Y'9�6�kj��=�ny(�xd���E�C}$��=�TK�45��pe���)�#m7�Zt��J��L�6睿�#x𯫑���sN?��:LP0Da�O�+�zc$���y���n
��SB���`׹5��K�0)�����h+�L��48q�$,\����5w.�JK�WXh���O�h���f[�0w�l�{�=���0�z����&~Ӧb��%(�<S&#3+�v��.�EA�v:�b;��O�&�h�J�g�����Jq�������O���	��T�Q���-�ݰ~+A���U���0�ù���`R�0.8�!WX-B�AksA�!�S�~�����ҨHl)�V�,_~>f̘�sM��������v���	յ�{�V�?�˖<��u��ƙ���&��NG^~�Z�i5i����H�Ђ����w󝽤���:�v/����5M���g����I�#��;w��Y�b���X� ���0�7�����8�X&�R#=�(p�ѹ�iy���\S�:OD4����6^���o�Tx���3�O%�S�"zG�E�O�~�5����I'��hr�T�����t2���-D$$贫kSS#Bv���|,���66�hr�+�0����C!m��d��sV��
���a������E����ä�S)�lE���ޛ1���{�r���d�R��IP>����َ^K[[;��F[K�/��°Z�蕟@���e���6S� k���� ���6���I��#���F��J�Uט���g� ��j8:l[�G����X~�1b9����h~+����ɸ��gP~ agu��ǙE�/����s�'��E[���H��1_Rי"�,Z��+6Z��+�~4i�!�&��+��b�
f%Q��i8}�y����c�abY9V��� �}p�]?��_��)�L�wu�R��o�ٹl��V9�^�Rǯ���@���� J�R�$��q ¤<����?�y��G>��/�g�X���I⼋.�e�\����
�)���M1� �Ӗa��i()�ǳ�>��_}͖�f��{>�~��]�Ʋ3�ByI9�M��3���k�v��;��I��o�~��t[�7�+m� ����ªU��5��'	D�p�����b�]#�� �V5�՗��pi7���>�"���J�#N�PV����7��p��[W�ʮ��J��q {�Vt`�����(ǦM��Sk����t���j/V�ơʽ<�V��w�����՞(�ؖ¡����I���?��I�����n[�+KLjZ�cW���T҇�c���q�Uf��'֬Es���zN	�C ���"7�T)�e��#�I���p��^F�p#1����͢��Btk~E�a����@X<J{<�>M��Td������3�aҤ��Vt�$�'�͡-}h(�����V�wl�=���t2���[ �(iD=�,l�tMm5�-���7b��}�Zn�B� L��3��IXq@K�vV�81,�/_����X�r�Y�+�=g/?�|�o�N�<�y��##-���(�9o�\lܰ��/���.=��A֯{�@A�]�O��#;��F[S����`Շ���QY�2G���ڴ�3�O&IA��2��-M�W��Ĭ�@� ��(�4���6��C?��$+����-�g����F'�u�-����mm]q�t�8��9	D(�d�@������������c'�5{�|��![ל:�Eq4壼��3qش���]��.��S�E �����Ix�6߾򬥈H<��c��{��n,?�t�M����^�����P�wk*@u����w�"�6*�������+� ���:,.J��(뭀Y��'����#�c�?��7l��o���-��u�l����vyc����[H_��xq�x��Ǳe��6�rc�����g���-�G@~h�^l۲�c�0R3sP6i*�n߆��Z������Q��U����O�S�Q���!�Q[�%]��l	z�+1o!�1���Q���n\x����e�KI�����f�kkkAue-��m
�6bc������O���ز�u���% N���Syy�(+-�ĉ�t���W֣֓!Ͳ�����fr�$!7+3g΅O�U	'D;�'�>H�IP�r� �H�!�<2�_y�ma�G���i��O'�'���Eb�y�d��^�
�_��`=��lL�'"4��9
$�1��bF��>5�m��_��5uM�iټys��m����
�Ɠ�@z���q����tn?[:z*��'q��ʤt$���1
O<r$ſ$�9�\ݨ�U���%��Ġ8c:�޲�- DD�G�ğ�xJ�7�ߺ��-���[%�5��K����i���_B��hό �|�0o�1�]�vb��}d��qp�c9��� �ӴOyY	�Bil�1ڲ`Eclo�@#I~!��
�J��o���ص}�1:d����Hᤨ������aΔ
Ȥ1M��],�9�Q@kzIew�q��������t��1��"�?U�I DIV$�ϏYs���{?���j^������D��Y�_��oN�����/�B{�x�������Ҏ�����H% ��zco�?k��w�\�D�qbȼ�C�G𔘌#��c��p��S@������������8��S�5�}| ����äY�0�������lØB{+��jq�6Ч
��6��W�[Ef�L�V�xKq>��j��)�I �7܀W^{���]ؼu3��ޅ͛6`�7��*�oތH��-F˭MMhlj���M���N�`�$��è��]m���Vt�6YTܺ�f��!��N���&6���d)�v+>� \!����t��1ҕ51�n��f9�s,��)���Q�)���a������
�hTBS�{��٧!3+E��3	>��,t��_���B�ۿ	}M�����׾*���ʱ�"dO�y��Z���8;]N�����Fmu�����n9���X`�}��<�!^ɉV�I|s|��'����AĘ��${�~ҪUk�_V�l��~4U����F�
Ǵ�[V��)0�����M��&��}W!���ib���	*�`����+�~3�o۶�8ph��}z����O��}򻪫�G3�������+�:;����Zm(eN�w�S�:�7X�H��[w���-��,'Y<-����q�өO
��TRt���r�m�'��3�-bys�0UOY�ɜC!'d�*mF84bGQ;-&�k��D�r:B���l޼ɴ�ǟX�g�~�<��Q(·��*4;s�H��Aښ������o��-�U�4.��r�
����{v�A]U�9�ˢ��0����d��)��!�ā�8 ���4��8n�v+���1��������_��W�d�)�n̚=זnn޴�������#�̉ӑ�쐅E\�+�����~�;q��F�,Yx*v�؃nmM>*MZ`� ���aX��a�f)�@$S��˶��R�%\t��t�At��&���͇[�ǡ������z�y�Qt6!��O�NҲ	(=!ly�5��Ǿ�vwN-���_|�	5 ��OQ�ʪ�O9,���`8�'����v��c���a�>��
Q
 ҙص��E�" �j�*�h����!S��=�c6��$&�>���Wj�ٷ&L���FQI	��܎���x�%%��t,?w%"��?�½��JK�l���C@�%�Q���3�-[�$o�M#V��3& �㽱A��!�4ף����d--��?b���q.�q����ʫ	"��g��<e��23r�q��&s�>io���z�S��XU[���Z�RT�g<@nv&��]D`���tQa��F4��&'9�Bd���Ӟ9Q<��%4�tb��3���T�����	��MS�n���"5ĺ�Bd���X�X$�����[�G�8�M��'���,].L�2�|�>l`A!�I7�6i�3m�}$����
J��}���v���ʷ�fk����������aU�m)�!*_��p�"(��ge�~TW������>_�6�QG{�n��ഷ5񜀇�zz��?�T�Y�!��u�fI�$�d~Y�T���
�Lo���"�Z���M�d��ttup�&PL
�/� ���|"�#b�#��W�]ڇ���Ң���ڂ��Fa��U��(���`��q鞹s���wh_�E���ǲ��1{�\j�1�kr���U���\���"	&1)y��a����硰�)� ҝ���lև�a�i�^�R<�O	F�|�͔�Ď�U�4L�2�"v�Sp��К�D�)�#�"fz4�s��	.���^q�ո��+QL�ZXPB�n��g�~���JO�^2,����I�2k5R-I��E�YF�}���}��f#�2�@GA�Bɯ��3��L�*���@%�I�F��%pim����6`Ӻ�h��BOW�\@�a}�헴1ƾӧ�b(2�A��e�h�0�v�����Dޗ���3�:�,!��Oä�ȰV�PPS{W�١g�� ��A�m�|�t�N�
��>1xѿ�zd1b��Ǉ헝��R�����M����N�C�8��Uv�g��PO/<��a�|'�� �� �#�|)b�|��a���q�҉����rh:��� �zX�䵗��K���Tm_pх���4�q��5�EeHO�A ���t}�#-5�m��7�^qrX'ъ��b�x8��2�� �Ӗ����|;C�A�m4�$���O��C�Q�9��o����	~�3ˑ�=QO��I� �a�C���1dL��\������p�����f�}Tqg��D�)A��(y�Me��X��"?������ߍ���hl�%�k �h0`P_[���C��Uh����JTL���C{	64���{�`>�������dh�VW�Q�<��������TW�;�	^���cG]M5�F}�~c9��V�Y�WWW� A΁�l���uzZ&���ŕ	�����dzK���EĆ�ŉ����sSh6�j�ZE"�����B����}�@BO
��h�S�4İ�tD�x�)1`�m
ސ��m��}��kV0&�Ӣ��ׯGII)�҇Ҳ2�O���õX��Ӧm�6���b�]�-��%���H��(����⎯݉�}�X�d)\�.;g._�j���2w�D�����_���O$c{��6�[��idf�b��������>twu���F�hw���J�-Q�1���+�ZjY��X��x /��2������@Ml��!\Ҙ��[�I�J[�'˱Oq5؆�;��U%���~�.��Jq�W��u�C4!�<::̼($�ö�BV.BN҈bw) ^mM�h%�<)��;Ʉ�ۅ
{9#F��H" 2[��j��kJ�E-Z�*�7��=&�y�Hôy�����m�&��w��}��+��,ljk�*S���m�/�& t;�z��H�
�7a�Mܬ���R��PQ1&L���;�����Ji��'Kb��y�
>?���?G �c"Z�|�do4E��P����Wj�&��1	�ǆ��b��2�f�Fbl��٧�DG[fϞeS�#l��!O�3;	D�:s��'�OGl������E��\ $;���XjZ^�P�iJ��G@��u�	��
s	��M�8�s�4��'��2b7�v��F�"��(ȔEP����g�ǡ�&�rJ˞w`�CHf^���D�:&9߃��v靖��G���A���y�����&g�m�Z�M�����.���.Z�X��Me�8�o��c����� 2���}��yţ@�֧V�h3�Ah3˞�.�.���:ğ��/�7����==��k"�i  ��a�-- h�R�������D�Ӏ�C�prR��l���=�ڇ}�y�݇�;wa떭��c���x�ŗ	��PT\�<�b����L�;����-D�M�F)��9�9�)(����V9}564��$s���_�H��h�g>��db~J�Ø4"	��ϑ�qA3�A_^�A�c�b�_��+�����.Z�&NĔ�Ӱ�`%�p���K�i�T[�+�Y�$GЊɓ���_����;�IF\�o?��W��W�Ǽ�����z����
�����K�z�%��.P�z�����<tM��6��OB���y�/hmn6����6k ���/��n��(uK�m���\������A�� ���/�,i����X|�r�7Bi���?�+���y�۾4��ԔC!D����"����1�e�����E�⩵�`���P\���.��(*)�)����������S$0*��D�I���H7yŅXu�*�~��8k�J���2L�:� ���=E���4�fk�(�%Mxɦd�\�Um�^����[�h��H�"24��:�;;G;�K��t�������3%�ܫ)DѬhY�:�&�X�i�%-�N5���r�ٵ��|>A��d�P�>k�J�	l^X��q �XD�【�W#iJ#%��b��E��E�k�'�0��Gp ��۝صsB�;(�:z��!+f?::{��W�ԥgQ�_����ޛ �uTg������}�$�vY�e[��;f� �d�$���$���%d#B62$@��	Y�vl0Ķ�o�%k�{Q��o_��;�n��V�,ےۭ>_�t�Kݪ�u�|u�ԩ� "@ݿ���0�4wJSc�T ��x-�|Sc�o�����Xc:BY!�(j� ���1�������k6IeU��7�4��h p��Ɠ�w.���
��o|W �j�x�:�E:%�F%"���ɢ3����LIUGV�v���7.��S����È
d�z��s$"�C���i�XLj��ֶ6�Z�5d����0�6��k�Sw���79�.����T��{bt;�c)ԅ4��b��D:�.�5p�(ړ����	C�R+���M�n�	%���`��P��P~�=��� ����[i��Yj�h<�}�Ҹ��TGG'ڻ::(
�hX�v���'B�Ә�����Y������{�U1|)�ؘ�ǔJ%���dC��:�L���1n���M���/��"~�ufe=
�,y��G��K�G㈢(�����|W���Ƀ?�1z�����+G�H\��2h�DKcz��r�׿#?��?/����KϺ�G�_}�2��5/�����B�0{a�cC���D�A��⛁�l�<9�r�q�6��Qk�����S��O��h�� 4B��x�Tޫ�8�C��R�ũ��7%���\iA��jFp=�Bh���"+J@X�,>�C-���%o޲U�g���wKEM����!��;�-�m-����g�ge۫^!���e4��k��Or�O}J6l�*��z���}R~�w�H��淣�ݎ^.�}.�l��@8⁆4����������w�)��{ ��;�#���{����?�s���`4*�8�c�ui|M�b��萚�f��`�^�)UHg$.�|� DbUl�c��p{���U�8�+H�e}�L(j��1����c=Bѓ�P0yCX�nL��g|(w��"�8I��FeM��%:��-
�	}���a(
���6.�J�\Q* �YˆG#r�LR��BFR�9x�8��<�ԓ�-��|����'_����kw���Q�Qh| �fԓ*R�G1�|�H�l8,$�M-��3�KKmEA��A�*j�2>��I;��� ̃\�H�+��x,�}�z��A�R~	���!�h?rx�l����7#� V(�(�ii�Ln�a\*��So�(ox㫤���܀���}I��4Wl3X��W���!�Ðq�`,�d/"�lU��X�L�Q��B���.]��4��Ieu�TUW�և��qa6B�A~QL�0jE1%���8�/����2��)�4����t�$W��̀�dQ�r�C9� *�¸H�H'��1�a��F�Fo$�AX"���xo -�� �oe�:�GȌ��� H��gA�[k��ʀ�ʈu�p��Ԉ��Rs�)al|���C�,�E#�C#��Tw�)U�	�9
d���ȖǩU�>["2|6�$�v\u��Eك���Y:�&y��_��H?W ����!��8)���}�<I��iC�&g��zq��������[�q8�׿Dfi��۶HKK�<�i�n�!���x�t�7��
��>bU���q��k�g�/{f��=^
?6�:����%�Yɡ{U����7˟`�lXY��9`�9⦪��$�i��Աx<X���fD�"�=�ø}3�쓍7�����=}�s���?�C�v�-�쳇di�"y�m����'e��{�;���/�1�����dEW��x�m��}����^�\n��V����o�]~���29yR������_�q��G��ZA7�v�����S����]�W_����ˉ�G���C~������Mo�5k�Kj��N~�Ij��$�r�k^%�\s��>~B��)�TU�MH�	�O�A�����]W�������'SRp&�3;���=,!~%��^c��ٳŁXe��u.���Nٳ�)��QG�YW�Է���Sz�{���VV2�aC�A�H�o���}>�P�Tu�(���d߉�_k���kD��F�{��Ųr�*ik�v��[�V�l�$o}�[��ox3��D��)��BI�2�U)��&��������dۖ뤣�I�-[�A�F�y�Z3�5-��s�惤��נ��ʐ��Ӕ3��@�J���˫ x+�v�%����>��@D5`�����/n����%.����;pd��z�a�^WA$��a{�w���ٱi�h�l�7�G��.�NTL��v�5Wɦ6��o�7p�lٲEI��-�d��������k7��&�'�p�]ј��뮖�7`�jY�b�rY�z��Z���Wɒ�KQv+@rV��ˤ�c�4�촵uJ[G�t�M��5�q�gn+�*A:"R]W-�ʸp��r	��*��(���TF%��8��q�l؀�Z���Nߩaa��Fl��� ��`v ��#+�3_�1���.��?A=.��ѫTU���C{��5�
Վl�i��d�TLl�
 lt7�
-=<tP{��V����o�o�Vi�G�8}����f(�L(	`��Au(S��jz�r&��7n����?�a],�фT㣆�V��o~���k��:����EN�8�U�$P��M�C����\�i|�<��c��/�4!p�������#�-ᨚ�Sm��Yv���q>ŋ�e����1��N��TS�@`˸x/z�4lE+�������_�� \���oC�d���J�m��(��OJ}e���/�G>���B�ڽG�鋟��� O��/��?���eI{���A������Z���� ���o���ʇ~�Cr��䣿�[��_�;ɠ7���x�������SG����vɷ��wi
G����cRۊF��0�7���ܗ�$��>(�!������_�����|N�A"WoX+�����=x��~��2:8�0��Ay� �Ay��p����O�{h���0�)��~�6Pgj;eæe붛�_�;9��r☷ �WC���o}X��I������w@�x�\�%C��� 	$��@D���-�Cjּ[
M�{hX�RٰxT~�7�Ⱥ��� ���ާ����l��(ǘ�9sV��
���HO��`z_%e�b����Z�|i��'e���������~<)GO�/���Ե�����M�_%7m}�,�;��CQ�
~� ��_~�.߹w@b�^/�����7�<#���ai�7�^�ݩ>)�g�uy�����������O���'�rĎ�\�]��9�T���+&wt.���*�	mJr���p�g:*�x�O�[��V�M���=�`8���_m�|�JK����}s��;�e��YGt�?�W�1!<GP�j��EҶ�Z6^�z��@�x�YjMٞQ�K[&�k��t�H�j��C�YjS��������x��Y1"�PpEjD(\�(������F�d�lؖv����zdDWz�f`��I�5��{�rz&{|���#��*�h *J=������g��j@\����&��1[��}�(k����Z#ЎL���>I�ez�O��#{�Ӿ���;e��O�>,�w�B*'��3��CKl �����aTذGГ��K{2i��!�}�'��Ɛ4���~��Ec�W��1�����7�I��<OB{
���PB-�E/�4��6�$g��X�+�~/���n�G6�|�l�^��7���G�yv^�j�t4�����?�qy�m��ukW��]O��g�!�|��Q��@������
��g�Y��O��<��#�^+\�tz�[�nUb_������J��x���ʟ��5��ګ���ȊE��[�(�����w��r�ʵ�mۍ�OwM�O���7H]U��ܳO��^�(.����,w�w�n9q��ј��)��u�v\�CPV,�e~�$�,SI�+1�u����� ���B!�7�%�a7���j���2�ߧ��Z�s�[�4�յ�r��q9���3��.*-�;WVV���sY��6��2V�Jr4+�q��d�zY��O iFO�B,�:@b_W_��@o�Y�ꤲ�Z+�+��4��$�X�<`�3w�*���FFǆ�Q�G~D��u6�nW@�oX�Y��:QO���Җ��GLpA>�5_H}�yjo���6ȸ�Q��
�d}2�ӧe^Ȃ$�\��EY�> ���]����}?|@;>�$�n&�\�����0V��AB2���[n�����䡇��֬�!��8:4	�ڝ�m��H�5Y@P^(-����刾�"��>Qԡ-�-�������e0�E��ӯ
�
���p�D#q�&MM)gUū�n���nFG��Y��[հ���E�ZQ�;U��ֶH�*틺��c�,�\!�-�Q�(�Ҫ�B@�k�������A4l|ـS��������eۍ7ˢEK  !�(PH�+��)a�F�];k_��.���~����s2�".oe_�F���0xD�(���Ɖ ���^������n����?~@��&���/�g������=r�������zB��1�\�DNی����e+dݵ�����K�H��T�OB�T54�Z�!��F�����U�A��һ'{�����GO��o�,]�T}��5.
ˆ��LIC(�w��@���#~��9�e�������
.S�����$�fC��l�O�3 
�)���cO�9

ל�)<7��hA�c5u �~9}�����L� ��Q�����������oC~�O_�Wy�G��&s��YS��c����m����K��+w��Ԡ�y�����'�R���Q�"��=�Y�բ<{�������^ee͞wRCLJ��i��:��k���6",S�#��%�%X�]����@}��I|�����!$�e��3x��}<+;w�Ty睯��s��;O#F�A�h��$��Ύ�@ĳ�
�Jy䱣��61<�
�5�n�/�G�j�z�j&\��cH��(�o�/�%�m9@�P>�������|���_���ݿO������:��&��)�莂qNS��P�C@��R�T��Ϗ�|�>��'hL]�
8�<d��� �J�O��:��۵��*oT�>�JЎ��mCC�#" $��֬^#�mm���y�+_)�~�+!țqHi1���p��ҩ�y�����,P
�_
l�&��|�El�ϕ�ŏ�����{@(�e�g+L��L�p�q6��k������a!�
�#���_����@hL��`uU����bRgϢG�FB�W;��>`���ϊ��}�PՌl�ٓ'����z�Ǧ����G!��4�� ����A����!S�����;����d������V5���J��|D6]w����T<�hWa�MM��iD�����&�������?���w��]�hI�<��� \��u-�7��-2�HIy�K�Tb�b���/���s�N-�x%��a�e۶m�ёZ��������:o���a��_��z�/_�ǚ��G|Cc���ZHs~���{yW��<�������w㶛��|�?-{��7�����ʿ~M���7�%��Z!l@�:�r};��Y�fy��'���^n�t�l�r#c���퓇�o��_�
�v9q�[>�?	��#�x�lٴE��69y��Ƈ>(?��w��\��B�Q�n�z������u��ǟ��zR��_~eW�놥��YΞ9#��}�9U4+@
w�=���j=�v�������p�+Q��7C���$(��hh ��j%G�����=����-�m�Nuv�ӏ?*cCț��!:>��i��� �+�.�]Ke�3;�sq���j�ƙi���Je�j��j�$����8*w޺V�b�8P#X.(�|��.e���hJ����������(g
-���X7 ��\�{8$;w<�35
���R�����@v�@:��VJg�rT��#��6
���`��wd��)���.�O������7�����	��\�/�����mm��3*��Y0N/~����c�_!�c�%���s�bY9���.Z�2Ƀޯ�a-��uU�Dlh�_m=�޸u�m���Lwi�rҲr��y�ǖkb�F�z������by��|V�@�C��٥6p���a>�Mf�[��k�=��ϰPp��3%#�
�f
�Zr
D~?G���1����H����1�c Aఋ�B�RC@����@����J�Z'u�~�܆#T�V��ǇA�M�^�0���7��M��*K��-7����r��PB�ԬN��=��I���Q2��0&�y���k�����G$��f��y����w�~��o}H��/�������'�T=�e����߃�Se�C#�(�-�͛6����A�u믖׼�5��T�-Z�H .o��W@�-������ ��
����r�n
5�[�k�pὼ
(
%-?��+�R��|a�.���5�`�����_��:A[��j��9'�ſ���Y��S���G�)�<��l�~��+*���V�9!\���M%���~j�N�e߸m�t.��E���_.y�E݀p�Z�R��n���{H���� �#R�%%96,��*Y�]UU+ǎ�����_Im}�܂w��o�+?��?e��:��0O:����9r��jeh����,���e�Qvw�����W��<������ep�D��A���F���d�-����C�Hz��3O?)�����_>���tpup��F�E��5'�h �xomn�p *9�у s�$�L�w����ť��x��J6�"�,��xeH�d��ċ���BV� ��bZNB��#�>��|����W���rߏ~$g�t�k_�Z����a���=y_Zv��Ne K©��B-'��7���!˺ւ�U"���P�4��Sغh'�~�����\$�W4Ime@�=q@
��2�3���bR�Q)p�p(!��C�e}3��A�utD��GR�f
u=^])� tI�v�:�����y��QOn�29��Hum�0&;v<)}�D�^u���(�϶�˃��q�\����jZ,���b"�J�qiY��R:PvA��h���v/>Â���	�G���J����Է,s��A#06�<�l-� �Uc�v������>��C{��y:cU�C��	}�6�.����gy��}�T�S��GZ�$V�e+V�Ï<"����&?��Up�>e ��|�_d B�=GB�ik��0���ƀ���7��-��cO�G~�#��{��X'�����{�7�y�,im�}x�7��m	'����3r�m����K�ȍ����ؤ���~��ݲ���;���|�ߔ�>���Iy�����]��������>*�g��L�7�Cj�] ���2d	�h�R��"�Q�2�{v�o}��r��)�����˽�ܣ �ٔ�=sZ~�����~oO��ݳW�~�I\��<���%r����C(�}ĪE>��ߒ�k�{Ƴ>��Oʓ�?�w�z� Y�>�-{v�{���t�9���fC��ڱK���/{��)_��t����l����~({��t�ȡ=��� 5�DǸ��]��\�v���Ꟑ�����ۅK��;����H(qc�� g�i�	I)5*M����x���o�5kր�u��5���Y[��g�&��Y�44����:�^��NA�Z�^�^�NFGF�4=�❑Q�T��/\)����~�$��d�JI�f���vY�Ӿ/�^25���ك'd߮�����\+���Y~�'�&7�|�`}�$�*�\�^��׾�U���3�2:6��О	���2ʥ��B|#�M�Nqi�
w�]v@��\W#�����هoD��G�b�Ju����i@n��Ab�H_�ڪ<t�hlQZh&hU[[�3���:@~��4��u����pw��N֭_����ؠ������]�����j�Űμ��L�:n/m{X�S�\(�\ʸ�ӿ���*�lA���Zy��^/W�Z����=����'n��&᠆C{�	���~eU���0���Zh�<�9h�/���l�ٻMi�FC���"=���~M�����'����3���|�C�5I~����a#�dn���F��R􉁰��gЛ�#��=��*�_���ɗ��%��'�DB��C˄����&���������;��v���k���Yѣ˛9]u���;vL6m�$u�ur`?z� m���w������W�
���Y,s�w�������L �i����d�$�M�At�����MH$X����e��Kb�_⑀����|��w�W��r��>�~��w�!_�����c���y��/~�o�G ��4Ȁ�؄!,��{��Oݣ��� �@�2 	G<+����/}�sr��'%3�/�H�އ~,#'K��<u�����'~�'��N�ɤ��#��Y/�z�;T�õX��P�8��h��r8""�2��$M�ʕ���������Q[@�Q�T�!0��>�e�	gx�D�'둃���]���7���@��#.~���y;!��%��:�u>��AI����7ʞ��N���u!��|Z��ů��_��<2��P%�����;���7��e�-��)�7�HF�s��G��C'A؎ʎ�{Q��Kߦ�q!���g�p���:,�@!(� 0� D�� ��;�xང�IsFS�$���JRx��K:���p�X�'���Tѓnw�Y�(���6Y�j�>�O{�a���%]]�N�?�z	r�wEې4��O?}�ab��	���VW�E���}��7����9�妛Ux656�G�P]��Ɲ���ؒc�
��s��k8D�����aC�{��P2�ڸ�"�8A�kѸ���@�κ�v������!����O���D���}{�8�lF_(~����Y�4Q��K�+�S~��.����#+�^#�����rB|1I5�Η8��4�J�Xx�����SOi�n�w��-[�n���j�J��|�&Y�|�pf W�ݳg������R��dY,�dХU{u�0	�@����8� z��Bi�V+22�6i��I�K�Gq���ĸT}R�H���j�,j���mrՊ%�4z�o����_x�|�ӟ���s�3y�R��:���/�tB�s��u�N�"��@ilI���0z���D�67��[�,�4�S7��ׅ�²`Ӷ�گ�Gɡ# ��P&Y�����1ˈ�n���*�4�,W�liB�\#�_��,WT��P���,�D���칶Q6/��C���~�k�p&���f�9-XI�+�����d�{�4Vr�M�o\����O��9$��*O=�S���>%Ǟ=)��_^{�+�w?����|��Z�B���擎9�u"��餮" �P��՘<��PY�%�:$^	��o*_��e�xJ�� �mr�9���h�9���jEF*�2�J�f�����0<�RC�}C����jv^8\96>����+�헽{w��tN��,��gcS��<uTz�~9u���*+Թ^Ck������p���`�p���-��p�F_*UɴC�߈�k�����>�4Ȭ��FA�ユ�] ��??Z��C+�&(<ؐsl�3ux�tx��Q0��qPa�����gEA�Ǝ*�]-�����u��i ���R2�5��<?8%9�F�ڵWɯ��}�����TŪ�o��3�iI�����KF]��$��^=1����}�x�� H�}�ݧC[�u�p�ȦO�;:dÆ2
r��Ӄ^yJ��	m�q��%,7�|��c��2^p�\p�v2�t��^�5�� 9C�I,J�W��@��l�"=����xD�B�X�X֬Z*�]s�tu�Bx��{w�p�p=Iן	�<���~A��~GENd#$"a��/�,�T*��=>j�@�4p
iDz9;9A�w��~�]�S�!����?��?V�V��z����儓33x?�J�Cc:+�������������z{�c�6u�ҍ��O>._����_�]s�l��	WVs����D'�g�v��(lR�o&:�:�W���U�'�]R9�C�e�ڤ�-*�_+��ȇ?��u�6Y��K��x�q�$�cA�Rѯ��F��<ZEP6n^+o{�]����ݯ�Υ�j�A�7���dOg��]������}u���^j�j���Z�-��j�<��#:���B����70$۷?��~�T+18أZ���JY��!�u����~A{�i���6eϾ]��?���o�+�������R[�P�#��ƔRk0�'�%_pp�`�f�uKK���O����wɍ[o���64�n�Zm�����f4N��c:4:��m	{<t���3Xu�s�*�PP-��F���W0Q�E����F\��XQU)���&!�sB$7���	+�)��$7������A�!p�?j!�{e��g!�A:�YI��%��e�V�����+V���m����=�^�w��]�� ���O_+I�%�pF�'�r���3ذ���Iy��ǄN��!���:	�#�($�Z+
�r�}���̫;���G�;W'q|?A�qŊ��I��#���B�L).�֭�5kVH%HgsS�4���ƍ��ګV�Є����2;���+�C5 �� m��>�B�C}��BN28O�� �
z�yd,�*�0�Gd�XR�na���Qx�~y�ك�t�r�q��5��Zѧ� ^�!��zUU]������ȯ������?U������;vi�W��M��A�X>�_�'AYJ�T�t��^9v�l�w�3�}�l��F\M��n�B aI=~B�A�cj!+d�/'�#5�������~����m����g���;r˫n�������%����e�TDk�~,R��p9~��u�u%�4A�l�Z�@�(gI錙d
u��fs�.4����^WS���&�t�]� � ��u\�2����� ����4ʬw�=~P��ى�ЉA]W�CH�hr�Kq�u-mQ���N ����9s��1\�������:%�� ��|X5 �2�&���f�:	
E(��@0� Z�z�W����N]���4�P_�x(��A���9�ī����$�h��c�<��"HPp�+���q�)����zz�P ����r>>	��J.\��i^H�h�O�D�h�OUnck�����ɽ���|���/��#�l�r��/}=�䃿���']��"�O��C{w��G�JGg����;gR�?wN������+TP�ݳG��}�Y�r��C�ڵ�KN;!7��ہr���_����%ј���,t�*�$ʞ3�<x�n��%��;A9�;�֊��^Uz7����=*Y�3����i��w�w�Ojkke���ء�eddD5�#����&��'!���G����dC�a� � "����9�u4��#p��3�xF�YT��-:t�+��g��!�N�!���a��R%*�����u�u�v8�n���s�L�桻�G��n�L9���vq�xH�##H���	{��$��q������zu�w��Y�)G%���͌J6��U��� b�U�.�%�A���N�+n].�HX�!�WNg�P�Ң��Ԓ4�� }��9�)\z5����8H�WQ>=�f�266���AB8�((�dA��W�����d�
xE�����[dP�i����=r��=!š6�'A�aA�'�	�ai\���$5tR�x�AٵcH2bC�Pm��\1#55q�}F?EC���v����dp�O	zcK����8H�|W�-F�鿃hր�l�H�X�P ����0��y�P0� ��Px=��P:Y52�U����*�6Z�@(�i3��#%�E��#0B9�]�slh���T!H���t� y ���Q )����GB\^��^{@���Ƈ�Z�S�S��#�t!a 08�PT�V\��,=O>��.Ž{�^9x�z�Y���EK)z艧䩧��S�j6X�l������ӧ��w�歲d�ٵs�.�=84,�=���Ԏ"�]�v������͛!6+���,����9�E�F�HmƤ��q~kɬ!�&��S� /[K���A8�P�wSs�t-[�Q�?��R�ٱC	��o��?F�>�hI������}q�%
]˜S!qo��V��P!�i�f�	������}C�j��ڀ;��R�ROO����A1g�d34rvCXJ�l����/�uydx�dPzA0{�{�Q�m'XG���4LF5���L�!5rgO���}4�\*�����6��뮓�7�,�^�E�ݺM��y���n4����s)I����%7�����������C"���8H,��"���G�ʘ�����WW/Xf�v���]��x���ԥ�����H2�C]]+k�^�TY��� ��ֱA��_D��/�%��]h� Hp(����K(�6T+��&)ֶJ!�#��v>�yC����C�����)����#lC
��44ԩ�w&���yBv��r���&y���"ڦxSp�VA�a��
\kfv��G�}!��'	`�#��v��%?�я���ȱ��[ϩS� $]���Ɯ����C�����	W@E�lĳ)��P��?���	�9��!��u���S��k�?戯�i��%38G�B����g�B���Y�m�I�E� h��)��.?��p%=��԰���˙�e<�W�L �D���楾�F*�QUG����ti��8~B�q�fA�@&8�wq�-��Ǵ�%�Z^��茍����g�{{z5<������bޜtyU��%�߮�cJX6�k�-�u������O8���:���՘���N���� 1�_��_�5!��_Z�r��X�C@����Q+@���x�u��C�U<0L���x� �4���*=XG��T�W����VF륋��Z'/�J6q�y���S�"�a\Ԍ�����e��vO���]9�7�nR���K��-�|�����H'�@4� ��&ӒA^�aH\^��k���ݲ��n)�y� �HVV^� ����oZ"�|�ը�)�qX	ߌ[�$�'�+ �˨Z�ȣߟ�O}��'����d�	�QPR���0�O��������W�"\�;'��Y���e�]R��������~�^�^��:�gP��~���K*�R������_޲H��~Sm�W�����] �t�[�՚��s���6&MM�ӬK�S;6��'N���A(A�Kg�"���v! ������7��l0��aD� !�0g��2�hYO?z�h�kl�31h@A!W�`"��o��R�ڙ�$(t�����6�� &(��qC+\��*��ˀ���>��!�a���@�����W�Z�D೟���
K\����e�3!�D���FrdC�a���G�T�"Wb�iao��<
K���dI2卪0�|�tЖdtdĄ�I�g�z
�r輗u�|�J�Jy$��3X�S0�L=aš2
X«�z/ʂ$B��rVA�E� JQ�z�fY�|��t�MH_D��݋x} ����G���'n�8���A�9IތK?~k�@ RphB�KӋLj$5eH/5[���H �yf��p ʋ ����ˠ�KqA�3��L`�P�	��}>���T�l��4(���F�KfR]Q�j�|2!i�L�iK~KWH�n��:�D?H��JI�Ꚅ���r�O~������i��t��o�z&��2̐^��is��M9|t�Dc|���E������5k��7��]��{xnp�� :���5[�+�m�l����^��ԉZ��Ir����n٨\�bT��_�@�>����F���)ˏߙ��ڙH���bqm�c�g�Q��|R�b�J���vݧ}��}L�l�����\l ��&�삾�s28:";�ڡ�g�v��ӧe�e.k�\7����hjWh�!�K�
�����7���"�V�NI���"jR(l���x�N�\OVs�-	 ۱R���O-�d�ͣ����xƗ�@�Q�@�@ �Bh�ID�P-�8#�8*s.��ϠAN"�i��;��&�x�؛G����݌�;�[L�$#K�T��Ԡ�y!0.������b��g��<�6�T�sH�e��A�5/�HP-jE�B�"$H|?;w��ۉ�:[��	x��𝐈�PNO���G�cq���u��l�f��-��8���&
"G*P[��	a�C��y�B�� �p˜iT���X��]�����2Er�DDߞ�������A�U�P�A�3����x߀d��&���Bp�X�,��v�Yy�܏r9"<xNBx߱hJV�,�?�Q���)!��CW$3\�D��@p�u̛˗3�c��r���D�^�!j��@[��iem�	K{�*	���*z)���=d�Fɾ���??$���J>|�$C��J��V�I�����{oqD����e�����s������]  ���$�DD�%�S��IO��h)g�AD��N[K��w�~�z���%�Imm��-3�����ED^8(Ɯ�e�B�����/'���S'O�TV��;���l9{�j()�|J6���(I�ӐP�a�aD۝�TUW�]���P��Hp-m6�2~Q��,:<�-�:2=\ǅ�]Z6��N"�C0�j�C��uu�y*B��Hh]��Uх}5�D>y�
>���#���Nc_.JG"F�I���C�fk��<���K���,��#ql�9܀4 O�L��j;h��6�S���D�Z5������o��	�a�4ʹJ�лt���d��p �C-�{W��t�,v��_����!1��һay�VW*F��Z��Giy0�1K̻^��p�P��C}&H�K�����A<�͐�N�y��$��B�Q����ȕ�8�*���u��+��,�3F��1��|�|�T��0�dZ�/�qyw�.�
\�����������gƤp.'թ*	��~��J����?z�lٲT���O��D�:���
:�e9��I�r�� ��!�
���L��rGZh��DD���y�G�9�$��Qԥ"���O��O�/���x��\"����VI&��b6"#��RMih������'�YB�c:�>���t�,��rD���2��ye)2M8��u��עڎp��/|����܊:�:���1N���#"�ع�Bc	;��m	<
Zz9��( F>twN�@!FaC_�C#2!�1
؞�^���CCC�ÃCjd��"�tN/�T�16>�k�У"�?>,cc�h����+�RPr�,�j����{�l̩
f�H��MR�L%u�[r6�$C�Wm�..��2�Q:�P��7�S�X4�*�(9�,G (�@,H>PV�A��}���|���āi�T��kYO��	�p�6�7I�����>�n�YN1�8�����mz�pb��$	iV��Lk	2�-��K�����}V�+��z��y�ls�Z�ؑ8�0��3)���q����y��̢.�f�� � ~�I���Q������8�-⧝^�Y� >�LrH��/\ԎS���!��'�		��F%v�>�"	u=u�_��K��K�~��2�D�G1����z�Ļ�ɱC)�u�%�����-�W�?�f�f}�T���u��'I')b��%�-W�u)t���"E������pX�������5��q1�t�
D�D�|��}���y��^�B��K4^�7��w�2E���'j]���9��-9����˞PC	P�����6�O
�z��f��P-;L?�iQ�t�z�e�V������5HuM���7�����+��\4�4ghL�p�w���jc�������BC� h�IT�]V�E!��\���툭8����^:�"K&��G�a�!-	�҅F�Ư4��
1y��mџ�N�U���:��>�8{�\7#���N��9�g�dd����0g�(A1>^C�-�I��G����	��tBN�����J��tG*bH'��t���e�ŧ�Ox:��F/�q�^j.B�O�HI�z��u\�CB��Ft!�hy�H�'�}Gf�y.&W�u��e1����+��c��b`���䏄���W����i�̃�1�u߯Đ���O�kyp�I0�i�|���T�<Ѧ���"��
����(Y� �j�W��H�s���4z�qu�i��o��,�>Ŧ���}���J�e$� U�n���b�;>�8҄���	������,���n��ֈ��Ԧ�RM#���=�^����~2��t�J�_(�}�_�_�6̀��ct�ttݡ�-�
(l� ��"
��ң[B!��A������<���O��8羯���8�3�(����W�i�Щx/K�6��'�f�ڟ�+k��V��V��	�����`z���1��ey��d��+��,5����7sM�U8���)��\� ч6m�ʙ17WOO��T�yz�'��/��Iv�s$����=s^�
/񾣿�}���>�n|�	�ꦛ��'�Ͽ*M��em�v��4"��î�R��qd&�7�+�I�}w�M�Un��ן�a)s�SS��ڜU�;T���P��v|v�"m�E�,�ȯeZ;����"HA�f��3��/?P�k���d��v4T_��}��Q�\tb�8�F}rC��W����z=g�K���Rq��Ǒ�I����1���56��(�"�a�7�怩H��m�c��tu�\��/��S�a�UċE��B_�fLa��v#�5��{�����q���;��iE[��6��?ahL�}�2��������誉r�����ۏ�@tE�
�f�f//��ߙ{h�)R��@N:N�m����.�M�H*�+	��n���e���A%R�!.�zꥧ"��r�yT�?�h�S��W�>�TW�!$?�T��4��D�Μ�ڟ�5���Q�؝��>��u���;��S;�������L��iͭ��0����{�*J�d�K�
r�U1k�2�~�������|j�J��^��cm�����ﰆ�	��0-�X�l��-��6mK8)��.�J��f%��T��jp���ꝧ�S�Aw�v��uYV����b:��'s��$4T�cT.:*����u0E�Y�����,�C�V�S6�v���t���;���7w_%��{�z�
����vŜ}]L�m�T�������n]���K�V읩5�1�X����X��X�5�:�ah�(8�K��;w2Ĝ�����kSU�X��}A809�m�gw�H����F��X�t��8���j�q�+G�Eo���&�����k.���铝���I��3��4�C5S�;e�?�P��_;1����ϙ�G��n�9�"5m���ȯ!��%�T���T���[��פT-p����>m]��U^�Uu�<�>j��40n�=ƪ
p�_�s��nZ�+Y����ϡ�%�0���4��6*�X���p��k����-F9�O2�jh�~}b�F^�[Ka�rΫ�'n��x����|���W�q�����[o��U6��)`�*� Ǩ=f!����eeҕ)^�B#�,++wM��r�s\x�-$��}Wa?�\��g���f��qϔ7��B�|VH=�l��. �!Zn��;��&N�������|�Bc �����(yՅ�\�x�%���_aga�)Ǌ�/��T!���#)���{������I�.��Bx!�m�үo�-Kyo��T��=�í/i���-ʭ>PB��<:�t��S�1P�����Q��u	�k^�������1SѲ������&7�Gs�����沛��ͤ�n��c�{ٻWZå��R�ef_�!�P>N��I6�D��@�!w"IX�K�ֲ�����m���\�ࠍ7ۜ����s������r���iN�f���⢈�\h[�eQ��O�}�³}��4��Z�0�����k*b,6�
!n��~$�B��q��7����H�|����"��G���.��Pڍ�0��rl�fs]�9O֫���a�on�-��gj6>˜�=h�(&��K֒i����Fc��C�փ������ѝ�=δ�hr�t%A��q�]��Dtyx�o"A�D Z=͗P�֒�ja�G+�N�AF,���)������Tm'�E����|m��
�l��s�	��gw�Oˤ%)��Ṳ�7����n����ܥ~!�i��6=7IN�A�����.�rV�Tp?�b�Bc�<y}6I�K����:�l���������W��9/�Gy*��}x����\��eY^��	R�����~�<=�<{p5U�z�'2����pL�)����j_�nk$��^�ϻ�N�p=��o-��]>�q��Ȯ��I���*��n�i�n�Jg���E&�D*O��9A�BrY�*��0#I��H���93�[�S��Ic��IP�:�B�4��8�T^B���������jk�p^�^Oj����>���pe>Η�>��*���?�{���S����
4"��&���9��N�f֖�FSuHK�\bZ�e������'�O��ٖ���(�s��+�U9��l��U�[�v1�T�qr�F������,�뼰�����������P�ҳ�3Q� ӵ���	cd[��e�����N�,�f���U�������ǭI�g.��9��'e���U���|~���Ƥ��LWR FV���~�/�I$SGu>Ea��:iE$�xu[φ%pӑ�v�8kԕ��S<��R�/=��0�X>rf0�����]9P?�ZŴ��|����DN�ό�u���$|腻��@���td��[�����n���(��>::a\��B T���Oȣi0����	�-~6-UΫ8���aӇ����NVCy�D��7Z�Z�+���ܯT�g�.� ����1x,�\����!�Ϡ�I�7�X�0���
��[@�=���5u"z��W���h�����b�B�o�&щ�=��U:"TR�
3Y夌1��l��3*T�c�ӌ�~�-W;�Tq�r�����=05m��?Z]	�l����vu���r����WM ���V�A@�I�^t��^���	�a\�YGsZ)���P�v�4;��������vJDrd=���fXY���zm��z� O���⌞h�Vc%2}h����1h�V᪜�k��\� ��6j2����ք�l���"���I�J���m�C�.w���(8�e_r�ME�^a<���N/\�e[q4�m�]pb 0p}a!���E����
�P�*���HCE'�����u[�لMyH�9,8�D��\��#��f�c�~�����9�HJv���ne�.	;�RN�����,|^Ѧ!��#��Eϱ���ݞV�.ʑm�2)*�jvR0��(V=���,"NE���^��&"���/.�sm�V�;}�f�M��HaUE��I�JV��!��ul�ͳ�$�U����k����3e =�2��%K�-�
��qe��m}�9��#�m��2F1����Uk�������v�	K����>`LM=�0�a�Uj�w�	���oF�Yhqp���D�Ã�ߝ"�'�j9�����+��7�8�jT[�9C������i��=��@�K��Wq�x��a��Һ0��:�5X�Z	 �-rǑ���+6t��;[4H�K)"*�~~�A'��a��H���x�r�Ac�؄���=�4�������IA�i*��s'հOQ�!�2��:�@V��r�&�b|��GT���
������m�8��[�͞o� )�껃�_ה��ڦx�AƵ���Ɗ�z��q���ᚺs �6,��\�E�r�*��(��q�l:�/�oԮ�Q!#������?�䝭�ۤ�7<��%�N�HDmy�/+fɻm�}.>^k	p�K��\p�TXZ%����J�N�:�	�l��0�����2i������Wy^���*8��Y=n�i�(��^#=ט��L{wYD)�𽏈O���N.N:�\3�`_�o՘.��*,�7epQ��Z3xG��
��xl �$%�2�ѾYo�����b�������ٲ��i��Z�"i�o�;r��v�чar�o�y��S-i�e.�y���^��_5�?4�L>Qκ1��<^��̅4�aU���/������ܙ��7�Ơ�GZ�����Y�d2 ������X��	Z��Z�/����� t�M�5(+Cdk��!eL8�C�|�p|��2�PE�������|��vwj��{�KZecl�HZ� �����R����`�r�X�w5���DM��tm��o(����܉\�i� `5`P�$L�]BC0������<�£����q6���(G�G�DH�^6���ċ+���L\�9֙$?�Z�M�-9��v���/=d��=[A�e�A���0+*��m����O�T�c,���-�Sz8��&��p0}n*Pio�PɢQ��.<�f�;�� X��m&?�~(���쌺��~[�P�%-=9��Ӱ��N�9�
n�xь`z팄�1���HI'�$��Z���hz'E���*�����k�j�*�
�k��1NŘ��� ?tl-+9�K	���9�T|�c�+X��/It9�����T2�%�'� �LO5?����6+>Γ�����֮r�Y��uL��&�+�)p�|0
�2����,4��Ĝ��**�V����n� r'*��<�(���;�A�8P��`?���4�l٦�հ$�,�F-8ߏ�w��uR��<�K���P��&�P�J��Vl��A�I�'�5�?O�����tFv�gI�\Pʌm�m��ԗ�m�#a+��V'�g E������[+��f*v�-Ʃ�����0T���t�ͰLIPzU;���&��ì�x��_:Jo?;�b3�SH �׬�N�B�3�� �A2�������6(�1�&����������_�B�������3D���	������X�nq��<��m�W�xg���7]$�;����S@�qƗ��@����3�ks�$���6
Bh�|�@���\���J�_4���̴1��R�b|��=�S�3�ot�pҪ6�]L2��(G�#0��'�"�R�s���<�U��'�[�~�=�V�8�ބ��F���e��)Co���t���+$�����gLLL��E�l��};>�>�u�{�7`�vSm��ݟ��	�����N쒵�/�yi�-�+�.�t<!r�XKZ	YT����2�K�c��d�O=�~�F�C�:�U?9�&|�=[�j�K1��mF��K@K��2�P<�n��o/oN���t�����_8u�1���jQb��@ _w!ngf�>�Ӻ��`�Ha�-k���-�+s\��Dʅ��A�^
�#�
*��S�����qA��O=AC�:p+i��o�_G�Է�і�K^�5��y?�0HC���7�P�L@�k������xY'���45;��o��_��At5��nKV��P��S�^T���["#M�JE�ǫ@|(����Gy��{���IҾ��]��6=�Y�$��2?���ׁ�ˣ��U��s��Z��?�������D���%$V�Kɩ��w)�� C䯞߷C�_8p��{��~!b����0U���K9���~��'K���Z�9����$�M��ч��H�/4������U���֧T���W/�}�rL\=\ȵ
��*T��CJ{D���b��r��i9��[ū�����Gz�d����]O�n�6���%�I��C��>�/�1�0P��Ku0toy��v�4�5�|�n�e���OW��뿒�͟~�Jc.����d�3�76��\/e&H��w���Z�d�H^b�����5Z�����N�E�ÂYC�ؗ�m����J��Z���������V,��{�_nrO{!���&�Q�Ƌd�'m$���J�0���U�Ԑ������T�h�a��v���?4x�yNm��0���}.���������Evy�ծB=* Y%-�Z������� Y�*��Ӫ��2�1����]���y�kx_]N*�A�C��{B_}Q��-/�����)k�Bf�Y㌧���-۳C�o��&��8RΓ�G$h���S���%=����9����G޵&�&KF~��T�Ź4�{Y�E��<�h�2N�}���=�1ީ� ��l<��]�j³cz�O.�h��,�N7����o�.x+��'��l ����%�xK$_�"(����0K0���0�9lh��	�$H/�KX��<�J>.Q˪�z��������]�]����]�����~߽ϴ��L.����k�P�H%Ӹ����&��ҵ@?)eo]�N+�_s��+��,q�ˠ`cXY�B�������4~�����	�>Z�c�=p�S��	��i�op�Џ'����ӏ�?�|VK��o���I�}އ8^3S������?y�)����v	Jչuo�_2��;����,~�^�P��|A���l^T��?�|����) ��,���P�x�� T���jOJ# T�n�w�K[#�+i|�Z����e�~:#��.���.�6D뜫��;��8W�V)|��4��2t*թ,��W���+Yq۝���+fކ���:E����缾ך�C�+5���@�����xS"9�%��W\"�w;G�����*�_I����ζ�8�����,�I<�B���SVw�O%�\�K��&�U�8y���i�a/}�ϼ�7�,	��kQ�H�W|��FU��t�G�$�K�m(��^:Ï>L�3�s����V��b;�ݴr�Y7�l�z���Zͦ�%G��g�C��A��Bܲ<k_b�8ڏ�WZ���� v����4��E�b�O��ǳ��YÆ2��l���^J�	 ��F���f��1�����O��]e�������5?����^�������=^}�����pګ����uP���r_=T�[�U��ME��έ��h7��=�Y��Qy2ِ� 9��~g��)GۡKZ���NoMK��T��<&����ko��ɡ��ռȇ�i�D�����_��7XZ[��Km����l꒍5�� vZJj�F)�.��t�F*
8@S�n���V	�`����wD���pj)�Fb����:Fg}1u��k~��^qV����(�������F���+k2r�ax���Ǖ�1�����yʰʈ�О"Ɖ�It��0�+'�ͺ�D�8�ع�R_�ZS�	g�}�]Z%�~��U�B�
�'��ǎ�[������|g��G�bY�7����b����:TC	�93�_J�݃
�$U�gԿ�D�])�1�Ԝz���Vظ��%�@(*��U����Ջ#c�3��qp�-1����Ѷ��E�$=�2pvn����oL��)b4�vG�Bis��av;��||�VZKmm�%�G����Rt����}B�%�[��L�(�+��e0,$���(�v;��s���~5
����Ŗ<)'��i
�*jy�s��!k��!H��o�^W�]��uĸ���_�/�������3�����p���f߽A}���5�K�6��B��I  2	éq����n��h*h�N������VZ�>���]�,�3%��Y_ �0��yl"}�E5o��2��C����O08���?:W7}��3�L�Dk7h�(��&����	��oY�D@�_�O�e�|hju]�P�x�x���]U]�r�f,���p�^_��v����)4�j^cccce��B�3��fo�%է���"J_bPx?[�4+�1����}g�f]���yA�O]ޔG7�|�E�c�~�\`��[�����{��dU�g���5:�j^�ɖ��j���i��)��gʬvVwĤ0�������VVV��	a�'O���805'.`�6[�[jY��1;��U�����{,v�W��m�l9�ii�5I---z7o>i���ZL�#�P�3�0)�h�Bw�鉞�h�7͞l��q��n�Rշ�w*���D��TJ&��Z��-R���:T�}t�!�Z�gX���)����˃`�����u�����*0ƞ�MƋ��-��G�+�ok�!+/�ei��v��?V4�*���M|���ϑAl�kN�Y��s|&��:�]��$�/�.KQ���3m���ն��Fh8�/�[_�l}��p��B�r(���*C�^2"��u��t~F��VH��E~�*wk1Ϳ��H��nf�(2���5�ڊϲ�EHW�9�4MtϜƼ�]������^��d����$���܁��l�jȵ.5�O�>I��d��E�����?@��dV_��1w�,�����?�6�LK"���A�h�ϐm���^>Y.���򸫴4Yٷڗ�x8+��ŕ�/$VTT4=��������-O�ab¦�h_�%���wO�]������·���:��4J�|�d��B=m�����m�i��7��*���F`��ꍳu�߹�{�����Y�o!��B��7��F�(�q��qU�w��.�,�%S9-���U����EU�F�ړܗ�e"%T���h �IO��f:�Un���)|��`���PW��j3b���HI�r��j:�Po��S8_F�>�&���_��ge������P���l����=�p3�Jw�N��ÊVNβэCiii�������
U��њ�YYV��sr���MWэԒZ�\���Lkq�h8R�h̝�<�w֫h�C{�N�'�x������'�_���4X ��nzD���tΌW��'���-���_R
A�/\�ي¯_�.���[�k@n��5��Ѹ�� '� oD;�}�b�%�nZT�eC�$�ͷ�Vk#�Ċ!����9�6ު}�戾�g�,��)�<-�U��c�8�tr77�&�����>�/#��i)�[��Y�^ޮ뽕q%\�{���O_Lw�%�{1A.�Y�܄gj�[�����,���04�4T9��z��v|<z�2�6�/#�@����g;���ly��{���ܜr�b�t��SH�#BY�_M��sZ;IiZ�,Y���m��c�$�I���*�m��Qk{+��X)�[6�fnΐ�tCJ�'30�)C�Z�k��C�l���U؊'O���*�ڮ֯?�h�6K�Qt�k��԰�D��WTk�I+�B�1`�8�o���0n��JC��jX��>9�?��ZϿo�d���\ٟ(o��Wu�,MR��7C�c>��9��}%;�
S�ub���]����p���vR��;j�&6�/�}r��.{H����x�ظXQx0�+;��c�-^Q֩g-v]���h��F�{�Pf#ug�S!e
���K��7�꡼�U��,+�T���1����ݘ��o~J^G�S�z���/����>�����~��ﳵ������m���;na��W[�U��{�aTd9�):��7� �X�w	<����;�V��R�}E���ܧ��F�6 =�oq{��'e����V��2�8����'���ߖ��n��*��][�7��!��:�ڜQ%�ϫ��=.��=�C6
���Y��J��-U�"��b"�2����k'ǣ���B�r�z��^j|(�1�4�|��ṱ�na㭻��IJ�*������
ە_^�������j��Am+v����o�N���jB*���Ծ��T��vf��&Ei}��﬇'�'���K^��Xl�tn��1zB�,�c�3|
��^�;MuVw�N����c�|�!��$j�oqY�xS� t��K���금XB�O9��='�z-��31^K��2�Y\\�Y���|9$W9}���+R9(Υ*H��s+ӧ�����5�Q����8
�xN*B���uQ@�Y������(kO�<C�Rs�t2W�7�*<3�� �B�~i��]k�����м]����gz�]�J��:E��ţ�o1W�8jzU*�6����4 ��bm^�]�%��b���^�1��Ż������y��<����y�Q���F�7���h�i$��L������+^��ԗK7�{��k@Vb5yk���$Os��uu*_�ҥ�V�S�سq���K7l+-,�=�;�u،��.�"�+W��D��Gj��wͦee�q�������=u��2o������2L��]ؗ|�����ll\M�W�m_�.��,�wH�TR^-�a����cە0����K�A�I� s�D��:�n/�<v��-�F��|��f���A����3�7��� 3�l��٘�d��ɭ�B� ���������f�u=j�Ŷ���E�#�?�1�՝��FJ����y��?�2ۥ3N��5�
�x��ХX_�{�{�ؿ�=��"���*���ϧ~|y3���"�@�%Z�_��������_�hL��?�_�?O*Y�z'P	L�2�r�1��j�R����c7����0�/�꾿zD�؍�v�ov۾,��Ez�����?n_�Ǽ�����e�B��^}霨|4f!-/��[�s�$�j��8��{�k����'T�(!�qӾ��ӳ��=��B� �l����"�!߿77���x9��m��F���w�>L"p��H��z�3�����V���}�5T#��M�./eҠ333/NIϓ���ǈ�����&��?�+������d1��[sȎ�Վ�����V�c7�E&��'_����ң����ଖ��|�!����g�MMMy��Yte͞	�z�Ap\��J^ћۣ?�Ӌ��o=��~�f�;,~�3����Fm�`v?�̙c�.��ز���G4����}����[������G��wB{�Yh���Qۻuӄ�f  t�CC	�j�vš�zؚ5�����E9�:^{ɠ��4{�Қ[]��]�Lk�U+ad��ql�v��T�@f����贛�aC���P������c~  �pl��V5�r�WMe���Mf2�N-�oRE���d�?~v�o����7��]�ˊ�YK����� ���Y^8�3'ν����\�`.jq�P(6���/ˣ8�<.��H�V��%J�� ��2�lÞ���15x�w|U�X�E�pX���m���]������{�f�����zQG�7?=���F�]R̩ؖt�#a/B�s�n����<T4�)���)�����#��]�@���/�a��e��n!�j �8&
HK����F]��h+�F�e
;j��H��)9]B�j�+"�_m��wW��6Q�fԑW|3�=���CSCi������~zc~v���A�J~]Z��~o	�Օ�^(XR(Z؉=̿"C���w��^���J��^��xC�K*{c���m+�޲\�!�Wd1����y�Pĝ~/pU$�~�Oǝ����Vi1�i��ض�N	��tϲtE�\:q��;!6�OI���Ng���[zn1�`i3?��qc:^���Њ�.~�c�_'�'��}�W�7:�>��ë[]���n١r�$׹���Dq&���T�&�eh�����x ������7���@'�p�`���ލo���d�&�6�W��^C�GҊ������:,�J�_k�t����67"Ztk�P�L��rt�2|�P�>;+.���bU�z4�W���*!�[~�sn���.� �)e��~��O�|8�wB8�h���e�'�5WTuv:Pj6��5�(�>�Ţ.Ϳ��T�?�z�U	{.1C���䮔�����-w䚆B�J��WC�돫Z�طp��� 9/�K2��@IQ�8��s��?δ��|�B\=�0�*㒓�pe��t��� Y��#KE�>��hv�Y�gVk�sP�}���z�Q.q��o��UuJIaI�K~��`�t��+�"X|7㠯�����)2Mo�c��c��\1FvQ"����#x+�*t
�����Y�z�Ѭ��$��4Wi^�_=*�K�w�������
���Ż~s�}�L���vܾ��P�T:J�c+
=/�]�_��$R�aR�ғx2L ��������F�"W����g��ܙM���6zZ�OO6�>��̯�?r=aj�U�5:|�9<�a��/L�s��A�Q� Irp�����^�>�e0��䑩Q�î��Z5�l)R!c�Z��8�S�}l�aȟ]�+��J��|h��񵎼��'m�+�ِne�d�!��p�f�.j�H��!�8^��~LzX������-X�FZ���>�lg� !�n���V��]V]���ҝ�����}�o+LV���7��ġ25�C�ޒ$��<i�^}��'��"��k!��[/�T�ϢǄj�SX�
�CX�,��
E	B��ʦ8<�,:8��©T�4Z��9AKW�EcO�C����l�~m����
�ȵ�~�֋|��$q]�VΏ/֋��j�|��JU��d�����%a/(�uz=Ui���#��ކovFF�k�t^�ũZX󗮑<����z����e��oխA�PWہ���W��~!���&v����?##��{ztJ�L�6G�:��9T���B8uگ�|��S��J_/�]�K��-�x\<�s1�o��hd1��'�yY�P�1�'
P�1���f^�н�yl�},���9�Ϟy�C�v(�����%V��|'�Я�gwwG�߸.������ǵ۪�� RװR 9�:	�-�F%'_���G��6���~� r�H�$Ԅ���D����B
���3Zo�z�[�@zz�"�����h���V��z�]�UvF���HKH����|�qߖib溈�����Dr�p��T����\9b�j�d��"]����q֭D�p�t�'?��¶N��X��B���i�hS���'S$�Ƥ�W%2ŧO��4�4*���b�ۧ�I��}��/��/{LM[x�����h�US�Yg������5?0�BJ*�/����$�I��������p�����Z̌���i�]�B`Z�>�$?���&�;�Yǿ�:]��K����������B"��lMk���Ҍ=!~�B�j�ߺ�Z���齟��*�L�Irϊ�܌.���^���l�ZzFqe����}��`y�h��+���7��������6P��	'��Wu��������Ȣ��7H�ت�fsv�G �&�\$Z�	M��eo�a�c;�����{Cr�ur��z%ʣ��0*?
qp�����`�B�i\{��|]�����dn<Kw��!A>�gŠ/��pJN��e#�"L�_)YԠ�������ʧ]7�t�֏�e^���2�� ��c�e4�j�peTO�[��(��c]�UEE�Jl��
ff,f��gzr�F�����q�(��5B��%k�NP����<k�}��k1�ዾ!ZY�1�,@��0%EO:}��	�V8�~dN��$K"�5�̛��G-�������񩪯�������g��y�B�oV�>�� ��R�#�{MB��:U�1U��o���'Ԩ(��1�?�����T���˹$��䆁Rc��]�#�̩�:zAIU�/u�}��ʚ�<��D�W�(��׉�Dz,f��J�|ie<;W$/)��7�J���`q
8_T�(��t������<�"ָk������!Z��J���͇�E�[һ�ZV���۝C��D��fm_&�ɵR��|Z�`��.�Bg\��g�[��;yt{3N#�JLܫf_����2���t���	�L".m��3�,WM�[�,��x���`��l2��t�,�q���T{�%�^���<�����
(�WP�+-H�@�F�f*�0�&�L0'E����ʁ<�ɟǬ���v�nRއA:�*1`�=!E���l���u���Øy䴔��9��rw��y"UG�y&��þ�׉����%�0U���0�0�C�6f����+����n �����,p��8��7�ɭ��(����ck��$/�ț��Q��Z��n���`�F�2�*�j�$Y�dWqiN� 2��7�W�ouK�p���S~P�mf;�y��U��*�I��2~-o��J?QS�>���
h�1>y`�go_��V@[�5C;Hކ)L�3�>��J 4dC��>���|�KG����F�g?��ُ5x�eƫz.�v9>�!׾m�J��k��a�aL{f���������a�}4�3Eh���&yY�������4�(�f�ry2
�b�<���g�4nX�L�0�P֔�~~��/[��#4?���9���Z���Я�f�~��)Ly�U��ޔ�!l�YG�(��G���sw9\���>f!�4�A�d}5��&��}�Эl�4+/xR��8�r�f_CP'���u'���m�EH�gNm�A�����-�ǲ=f'�N`)c�H�
-	�Gc�X(*v�X�S��P��u����AC�w'xD(5ZT@J�ђ�8�)�2`�>���L��Iݓ�W9Իa��?{�W���G=�ȸHD�]�_��۶�0d��0!w	C���J��CA�ԑ���B+1a�;�(��^O9����-E���m醧l�*c��s�^����yb��қ��ͮ���%�%#`��ooC���@����~�Yi��-�]�%R�n`|	˅,)p4p�h�V̾���r��ۓx��+r���6#�N[v��O�h|S�;�|3����oU	ޒ�ݭxz����ݲ��a��^H

�`��*Ǯ݈��EВpq�{�&����6��Jb>�x�3�/���Yߌ��{����脱K�,R`z%��s����;���J��oįGѓ�9�����*�[[�׾� Q���YV�G����<�n��I�Aj��L�.�m�ɗ�FkJ`����c/}%Y�H5q���ЈQ�R�͸'���4,�nf����>7�+?kO�&���Jl�C�t��L4��X']�8�d�`�t�.�0D����{� }ǫ~%8~c����i@��>��a��'k}\����Ѯx 3v�c�H9��;���>e$%�{�)�w�0��]
N�X��H}���4�b/a(8�lm��sݘ34�gc���1|w��m��o� %�y7nw�Ⱘ/B��6Z�._
�s;p��s�ݟ�$���a�� `����TK)�����ץ���-k�M
Ò@l.����^Rr��tOSϠS�
��θ<�D�#� �(�*<̾>����X������G�������8��"���b{?�\)���y��±8�4(]�ia��${�����Į�u�>�c��Ӥ��jҪi��b=3@�]�DfU��
ٲ%��й���mqr.��
,�-�7hN��X�,t�	����SXΘ)�~��ug�02$M���KMΑ��	��bI
$1��qy"'��^}���������&����+D����a>E�)аj�DQy�鵭� ��`�Y��S������2�Zuk��r3!�f�]�j�!���B3c����F�!��Iv､J|_��Q����A^.��(�x2>B���+�>�
��n(a�����zz��`�a%O8B� G[[�e��d%i��Οg�@���Œ�	�6(8oZ�]-���(��5�j%�aւ��n�t	��B�-1�!{H(n��Y5:����&��z�_z�xQm:W��n<�������J�6ޯYq�P�q��:�9�4L5O<%��f��ELcc�Q��/�I�'C��4�U�?F��|��6m���N}�Pa����(�����LG=��q��-XG�o[�N��z��"�FA��dݒ�_��sL!�V���z�gVˈ�(k�a��9�k`�x���ǟy�^p��P���|/<4K9�>�=R�c1qv/ӫ8�=� ��*a��T�����8�ݯ^�z�A������;x�0���ǡjT�E�N���w ��pH�T3����Y�P���4�D>P4�*�/�kU�־f�$d�1��QFF:xr�[�ףd$IgNϦw&aYq���<��n}*�t���Kx0��C��~}m(T�_�er~��AHB�s�r}��)��ya�����������KR�%�x�$#�B�B$#�NK�ݵ��m%�r��d����N����-B '\�SQP�ttR�b�\�����0�*�>LȠ!�˗������mB����`MY����I�=Zm9 2*��B��g�t�������/���3-��@���;\�4������"i!c,�/�BXh8@��_��M	��]5��7G+����$�Kx�A���M�w��R8݋�C�^�p��0¨��h�*��
7��G��pn��Y�PBr#C@R3� 7Y	�����ϟ��zf�i�Y������g�7�7h�1�� ��Iq!���l9�=c<=7�ܧ��2]����Ey��;pB�c.˭�"ill�=�\
,86|4�m��w�3�"���
�� I�v]��3���"�X���\֨�����8���	<2�@�Ao2�'�s����k����I�aT�L�� �� u�C���7
Z��w����q>纤E����2L�-����*�Aل���jc��������#�=��K�	{5lr��RU�^9�L�3����:��s_�0���Ґ���^�I��I��ʱu���KD�eފ�������������-�`�� �XXBTQ1�/�j��o���|�H6;4�Au��-c�g7%�}�rz/�`�㿟��8���$��a4�����|Iw(�P�'���j|�j�ԥY��N����`�'R��\�7�h���U���+�R�x��)��n����|n�|�a���<s	G�����{.�/_Q�������q�(���0ʓ��.��A��� ���_�JGK���N"��1�Q�1�� PK   ���Wl�#�;  �     jsons/user_defined.json���N�0�_��Xv�4un�^z �'T!'q�J�섪���J/P���3�f��w�d�ڽպ�k�O�<X�F���2H=)^�ǃ��ru�i����T�7��QE^y��F�#5j�,/u�Ә�s���XVI'��g��2�f�	qN֢w��	�оr��S�s�G�����l�ׁY�ƒ�@̰]��Z���-vHA3��������P�&�̲	1�c0�1`���z�������C�s&���RF���B�U�oM�n�OͶ���B��w:�Hg���k��%����>��y:�8��_�v��p<�p�5�\߸� PK
   ���WHX(�  Q�                   cirkitFile.jsonPK
   l��WK��( � /             C  images/967be514-0483-4001-9c2f-29bd6a1b95c6.pngPK
   ���Wl�#�;  �               � jsons/user_defined.jsonPK      �   (   